library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
package ramsize_pkg is
  constant c_lm32_ramsizes : natural := 458752;
end ramsize_pkg;
