// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:02 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bNZ/isRM7AY+Ok1iU4viU4A0UzIbFYqJyI+ebJyLAkpVD69Dn0GVN5vUnOPUyOec
xPYhIKiw3NQ/3MvLOBTQN3K9/PNuDhtSahsNANiUMD8ssfdJJPfBSEad62arm4XJ
eNayNkJ+rIiDWogQsct4bmxX6Stn6Odj9qNteKWREVw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
oPl8oekdwKD8te7CoeXEFIbLN6GUHQWOQ253O65EZDL4XrzzkXCv1mo1dh98inUr
8i9zrP0jT3qiR9tkb/d1IgzghIe6x4DU6dkL60HZN9TCneFFHXxdxy7b/o6oUlVX
o/ySttQ7bCkUix0qzElA+gXnukdF/WOqbLTaxA3Ab3GMgUQZEzv3MMAnzxm6i4xL
OkEpL6zRkIhUK6rlln+m+5Kh9ER+FYH6Vj/qMV5O36urYG4O2fsTqimfN2g4KIsI
55FzDDgH9reJZOr/86VmVOampphV9e47lEw8Fkzq98MmJbnCKqwLYZHnpTfIWd7F
zfC7Lj3xLLUxPfTB1WXSHUtwm1WnNcEkKhPhfPs6/qo9HdyRdf8niru0xEHQI20B
RQH83z/B/9dEo+pTwzV/JH6+2nhQy9uDesiCUwIA/nm58TriMDMh+3smPZIXCGrq
+84oOLV3Rh0Y4qI/nB1nYuNir+c0pBlnOz9ex6PxJLuAS3VZ5kcsHY7CYr7RjCXS
NECF7mwlSEWy9gycvUU3SD1RRmLX1IFyBKynBcne9I6H37sojiOOr3ZCCffKz+2D
4/o4nzP9DggTiPwiUKN3i2zV5llEJwGUXUUusnCBxGgNNg9tcgde/ew0hiBPQfxe
yjGFO32dry0aVvYeXCWml0ThWozhKy6ya82Xm480SxY3GY0GKe96ui91/7MvoTWE
Dg+iYrQm9ZPheIWjQOjVAgymm/atXJTDnim+vzPkrvIg6hg52cN4Z4819dTp0HO1
DBgYxFrJ7rjyif3Pm6G+yFOV33LYxe+QSDPY4bUu/guXPuf/CYskWJNKe0LOA5tl
m01O3yz4+YTN4Z37M0VviWejm9WAn1fDgT1ABwu8pmA3hyKT4Ylmp1ndP5UBVyzI
RlkglBgVjE6IF0c9wWp2Jz8cjvFr1ht+Zt7mTK6OC+BIC6N+TMm75frG1ud9nSZr
sXhlMYRjxGcTM2q1uwTIJtMLvuSW+2fU1CTRuKvp8C37TtR1v4JpZ0bIocJsyl8G
dyNZBZqCUoHinUvFqbSaJiWX6Gev8SC2tciL6vbuYR/mX0JWZj58yHaCyHjC8Cxx
VUBK2bRqR5wD5XGIREw7mmUdblaim9anV1yl+YVLoBpgsrVVVx/DeacYaj+CzKIy
/RPtuK36b4AyU0L51nBYBH3thgqJA2q6DJx32LDz8Cf7X8vmXw+olWCEctZn9ul9
GvQiY9/lrymopK6/UbrAbiKDLnjq4CBjozJ93wysUfxxFdO74Urc/QPv/9gfq7lU
qCjm6tqjpxg/kd/ky0LtNagiCfI3uvXprBG5NRNizW3ZJN/aztVXEfXn/knkQfi9
6IueGGEjJNThqZqWzfXfjQ71ZlCT6HOiawoSajag8yLPzJq75Bio7RuSKUbhtsZG
gf5byLrwmpw9fAxYfvAvJBR29aE7hSHu45icq17edAYx7DPJ3C53Dw5+F628iTAb
jr8y68T+v2Nor+xJRPobmbDWJcttwR++N4qgtrzzJ+ymZkKbhRyKKVD1/NNaZXuz
XN+QPEIPYY9HOA4kF+oamNp8JKRkWJpxxVgjuNN9VTfj5mJxHDKvyubmGg9jBJlA
eP/rP/j0ykPiOGpnOCKEuI6k+7j/tOZlXCRcl/UzBuqS9psb1Q+bY7/76UVT9ozN
+IE9+hnLY9zuptf0PiG9p4e1/eRwIJt8IOGKDrCn9ofguyXSR3vsJh1EY2AUs/a9
1WG81yMQyOf7pn1esu1H/1JEVictWz67S1aMKeTnoz8eXvriCHPZjyqCZoQU06cE
2OHx8s3fCSvQOxFSx0EMSvEASXeAh0BsAa2ZaRZEpT5cSmTnq+s9uD5jADUO/WyH
KBeCa0qjFAQKPXcrfjcqq67t3UcGU5knZvoLHgwFE1yee2rmMifp3gz4ZkaoTiRM
iuzN4AleLyeGtYldgrHvYwUx383G23SIoBz67PN3vv5vEbCOho/o6voUE9ksFvue
F66zz0f6K4uPZo5BWpHe54CjLWwjRYGzUVfEDj3fkwsbqWrF7Nf6QtKCm/m3KGdh
2Or15I8fzVyJllnv+UT+JfwRgjZZ+UkS6+VnlH04ZwUvaUwuvGbdbxZK+VP+4RXg
1dgoe79x8l8RU3HWOdDNtZKqvswY7tLxazIu6HhzLv2Tkd/O/naogPVpIqIeLgYx
a01hFHBdv2DN1AEuSM3zJqMLV1gor9A59io/PkxMtUgSBDW/X81oStkm7B2chAVm
+vrdu7paHcXg3DgO9DGm5fyLgwb1eiQYuBCgzWgwCqGit8wFuJLZgQGxAQAuiRc4
PWwZeYcGblQcX3GmpDjClI3oo/EDjhPRKw0xZLkWY/9542eOI7xFeD4QkadukfYX
xDV9ZNoO3M4tXlzWad9XFInBybWoESwxWLUbKT4/nURD5wuCu2a2VjavJhM13/SZ
1+as9d3Z1r1tNh9QEkWF9YaEQdIKK0PtSnC0gNTpNKcmFdpC3N3wfKxJGqorg+gY
G4THgfZvC5UROZ/Z4b2egihm4eZSgzUzrsIUEqT2IvaL0PDAP0fDfshmv1Muuiki
7DxKhl7ydTrEAtEmhc8fH5IUnYFBfzyOJMmIkSAY1ejSvMrSu2VSFWObD8o+TE3O
5XNfmquIhX/k5/W4VjWFmyc5sbbM86tyUG9zzlcnjnvWXmy7ybNDVOPSqcUyACvu
vODXvWYv/EyD/J8GuQm7v7uENREIA6NC6OiEsgFIbdN3WyEsIXhR3wzrBZhJlGhY
9G+aOAQ2/hj1/PBqZRbO5Gj3ce3Z5tlSTEbzSXMT+SVoXuMJEgTv/+ZwcJarje6a
yQzNZoreRwPiMiKj0WgqJngN0TgkD+55KT19Ix5pWQuydm/qU4SLISt2T7btvzhG
avpbI7fhrGyQsinkagbj9UwZG0E8V8kRE/KN4WFOEzKYMR1HOlZLw6zMFVJTQrh1
TTD8i0fjsZtvsz3sDbvyYRJIM1+0/zDZU+YZM6W5zoumPg/fNao2YFwxid0eM33R
rQ42gK2eUZBfPUJGkFi5i0xWwJhIGZkW5uJ0v5gGFofvMY68zS4gAICH/1YOjQ+s
9cNcjSWPrJR7tYF/B4sbbCoo6Odf6StUcrFhEZis0YrmYfYngUi1S0xD8Y7uhwqK
YrUM8J5xa1QwhmCrQrdeMY6+kHKI3Pk5lomcUtSTByd4pTWWvL1KtS7z+gc3KNz8
QXZjkJmVdiqiZMHsNY2d/MgCr+RSjuivITWFRu4Q79TattzdiwBUZGzoqOMu2prt
yx4MqOZYc3gcdivoXpWEG4MTyRKFJNh1p8CZj425NrRQN1rxByeN+EpN3xiDUztl
xr0HhK20EUjmTNTrSgZTJYeu/29S5GNCgdszs42dEhQ43TMXax4TEd+wyNp+sCRC
ubnQB9906TJsUohN4B1Ho50pWQk4DbaPVd4ef9kJCz9M/aaZoA/r4X9VdmIHL4sQ
l9rqLSl1SDBAIF1W48r4H6JW+Ocs41foEMETG2Pl2oSzhGyh/BJdQpLmB9U9yH8F
fXXouSet5K0KJi4ynzKwpipHYvyF0oOmxGnPpoq8Db0ANKnxGT/Ij542FKxrvWlZ
xI8ExJE6DsJ9kCKLgU3CcIIzmTvn1dE9utDK+9VzeSCCUfFe2FqXIrmkq1EG/gm3
XF5dyOxWcjZQma4R6+vh6o+KK1nzJd7PH7ll+Y4cN67pY4uZhAPp2lNOvVBBuIoO
XS2LiOE0Uw1LZx/dn+RuYd9DvNND6LetakL183FZI0N7lGYdBWz6KPLm8EGT0U27
d+Z99Scja/aB0qHx55EJC5TxWskoy0dq1RchgF2Oh2js4oIyrtE7O1z//WyKaTDz
HdFopemRpuPESfoDqZDjuSIhlrZC6Rk8tG1pyYUE8fQziJUddqJc1XT6rrvpOfvo
NgaXXxpXyV9d/BukKJ0U9tkhJhiMU9SJ099CnA2qPzBhzkByP5n21t9eNBeHzLhZ
fEIhQ+14piV7J0JFaLWeeQ==
`pragma protect end_protected
