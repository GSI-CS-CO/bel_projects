-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 9.1 Build 350 03/24/2010 Service Pack 2 SJ Full Version"
-- CREATED		"Thu Aug 26 16:54:14 2010"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY chopper_m1 IS 
GENERIC (CLK_in_Hz : INTEGER := 200000000;
		Loader_CLK_in_Hz : INTEGER := 150000000;
		LPM_Ein_ist_1 : INTEGER := 1;
		ST_160_Ein_ist_1 : INTEGER := 1;
		Test_Ein_ist_1 : INTEGER := 0
		);
	PORT
	(
		A_RDnWR :  IN  STD_LOGIC;
		A_nDS :  IN  STD_LOGIC;
		A_VG_K1_INP :  IN  STD_LOGIC;
		A_VG_K0_INP :  IN  STD_LOGIC;
		A_GR0_APK_ID :  IN  STD_LOGIC;
		A_GR0_16BIT :  IN  STD_LOGIC;
		A_VG_K3_INP :  IN  STD_LOGIC;
		A_VG_K2_INP :  IN  STD_LOGIC;
		A_GR1_APK_ID :  IN  STD_LOGIC;
		A_GR1_16BIT :  IN  STD_LOGIC;
		A_nMB_Reset :  IN  STD_LOGIC;
		A_K0D_SPG :  IN  STD_LOGIC;
		A_K0C_SPG :  IN  STD_LOGIC;
		A_K1D_SPG :  IN  STD_LOGIC;
		A_K1C_SPG :  IN  STD_LOGIC;
		A_K2D_SPG :  IN  STD_LOGIC;
		A_K2C_SPG :  IN  STD_LOGIC;
		A_K3D_SPG :  IN  STD_LOGIC;
		A_K3C_SPG :  IN  STD_LOGIC;
		F_TCXO_In :  IN  STD_LOGIC;
		CTRL_LOAD :  IN  STD_LOGIC;
		CTRL_RES :  IN  STD_LOGIC;
		Chopper_Clk :  IN  STD_LOGIC;
		A_I2C_SDA :  INOUT  STD_LOGIC;
		A_I2C_SCL :  INOUT  STD_LOGIC;
		A_AUX_CA :  INOUT  STD_LOGIC;
		A_AUX_CB :  INOUT  STD_LOGIC;
		A_A :  IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		A_AUX_A :  INOUT  STD_LOGIC_VECTOR(11 DOWNTO 0);
		A_AUX_B :  INOUT  STD_LOGIC_VECTOR(11 DOWNTO 0);
		A_AUX_C :  INOUT  STD_LOGIC_VECTOR(11 DOWNTO 0);
		A_Bus_IO :  INOUT  STD_LOGIC_VECTOR(5 DOWNTO 1);
		A_K0_D :  INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		A_K1_D :  INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		A_K2_D :  INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		A_K3_D :  INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		A_Mod_Data :  INOUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		A_nK0_CTRL :  INOUT  STD_LOGIC_VECTOR(2 DOWNTO 1);
		A_nK1_CTRL :  INOUT  STD_LOGIC_VECTOR(2 DOWNTO 1);
		A_nK2_CTRL :  INOUT  STD_LOGIC_VECTOR(2 DOWNTO 1);
		A_nK3_CTRL :  INOUT  STD_LOGIC_VECTOR(2 DOWNTO 1);
		A_Sub_Adr :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		A_Test :  INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		A_VG_A :  IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		A_VG_ID :  INOUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		A_VG_IO_Res :  INOUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		A_VG_K0_MOD :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		A_VG_K1_MOD :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		A_VG_K2_MOD :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		A_VG_K3_MOD :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		A_VG_Log_ID :  IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		Loader_DB :  INOUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		Loader_Misc :  INOUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		nSEL_LED_GRP :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		SEL_B :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		TP :  INOUT  STD_LOGIC_VECTOR(12 DOWNTO 1);
		nExt_Data_En :  OUT  STD_LOGIC;
		A_nDTACKA :  OUT  STD_LOGIC;
		A_nDTACKB :  OUT  STD_LOGIC;
		nMaster_Clk_ENA :  OUT  STD_LOGIC;
		nSlave_Clk_ENA :  OUT  STD_LOGIC;
		nIndepend_Clk_Ena :  OUT  STD_LOGIC;
		A_Master_Clk_Out :  OUT  STD_LOGIC;
		nPowerup_Led :  OUT  STD_LOGIC;
		nDT_Led :  OUT  STD_LOGIC;
		nSkal_OK_Led :  OUT  STD_LOGIC;
		nID_OK_Led :  OUT  STD_LOGIC;
		A_nK0_ID_EN :  OUT  STD_LOGIC;
		A_nK1_ID_EN :  OUT  STD_LOGIC;
		A_nK2_ID_EN :  OUT  STD_LOGIC;
		A_nK3_ID_EN :  OUT  STD_LOGIC;
		nK0_SWITCH_ENA :  OUT  STD_LOGIC;
		nK1_SWITCH_ENA :  OUT  STD_LOGIC;
		nK2_SWITCH_ENA :  OUT  STD_LOGIC;
		nK3_SWITCH_ENA :  OUT  STD_LOGIC;
		Loader_WRnRD :  OUT  STD_LOGIC;
		INIT_DONE :  OUT  STD_LOGIC;
		LOAD_OK :  OUT  STD_LOGIC;
		LOAD_ERROR :  OUT  STD_LOGIC;
		RELOAD :  OUT  STD_LOGIC;
		A_nGR0_ID_SEL :  OUT  STD_LOGIC;
		A_nGR1_ID_SEL :  OUT  STD_LOGIC;
		A_LA_CLK :  OUT  STD_LOGIC;
		A_nMANUAL_RES :  OUT  STD_LOGIC;
		A_nINTERLOCKA :  OUT  STD_LOGIC;
		A_nINTERLOCKB :  OUT  STD_LOGIC;
		A_nSRQA :  OUT  STD_LOGIC;
		A_nSRQB :  OUT  STD_LOGIC;
		A_nDRQB :  OUT  STD_LOGIC;
		A_nDRQA :  OUT  STD_LOGIC;
		RDnWR_Transceiver :  OUT  STD_LOGIC;
		nLED :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		nLED_Skal :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END chopper_m1;

ARCHITECTURE bdf_type OF chopper_m1 IS 

COMPONENT bus_io
GENERIC (I0_1_is_Input : INTEGER;
			I0_2_is_Input : INTEGER;
			I0_3_is_Input : INTEGER;
			I0_4_is_Input : INTEGER;
			I0_5_is_Input : INTEGER;
			ST_160_Pol : INTEGER
			);
	PORT(To_IO_5 : IN STD_LOGIC;
		 To_IO_4 : IN STD_LOGIC;
		 To_IO_3 : IN STD_LOGIC;
		 To_IO_2 : IN STD_LOGIC;
		 To_IO_1 : IN STD_LOGIC;
		 A_Bus_IO : INOUT STD_LOGIC_VECTOR(5 DOWNTO 1)
	);
END COMPONENT;

COMPONENT debounce_skal
GENERIC (Clk_in_Hz : INTEGER;
			DB_in_ns : INTEGER;
			Test : INTEGER
			);
	PORT(A_VG_K1_INP : IN STD_LOGIC;
		 A_VG_K0_INP : IN STD_LOGIC;
		 A_GR0_APK_ID : IN STD_LOGIC;
		 A_GR0_16BIT : IN STD_LOGIC;
		 A_VG_K3_INP : IN STD_LOGIC;
		 A_VG_K2_INP : IN STD_LOGIC;
		 A_GR1_APK_ID : IN STD_LOGIC;
		 A_GR1_16BIT : IN STD_LOGIC;
		 Latch_Inputs : IN STD_LOGIC;
		 Reset : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 A_VG_K0_MOD : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 A_VG_K1_MOD : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 A_VG_K2_MOD : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 A_VG_K3_MOD : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 Logic : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 DB_K1_INP : OUT STD_LOGIC;
		 DB_K0_INP : OUT STD_LOGIC;
		 DB_GR0_APK_ID : OUT STD_LOGIC;
		 DB_K3_INP : OUT STD_LOGIC;
		 DB_K2_INP : OUT STD_LOGIC;
		 DB_GR1_APK_ID : OUT STD_LOGIC;
		 DB_Valid : OUT STD_LOGIC;
		 DB_160_Skal : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 DB_Logic : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		 DB_Mod_Skal : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 K1_K0_Skal : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 K3_K2_Skal : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT apk_stecker_id_cntrl
GENERIC (Clk_in_Hz : INTEGER;
			K0_APK_ST_ID : INTEGER;
			K1_APK_ST_ID : INTEGER;
			K2_APK_ST_ID : INTEGER;
			K3_APK_ST_ID : INTEGER;
			ST_160_Pol : INTEGER;
			Use_LPM : INTEGER;
			Wait_in_ns : INTEGER
			);
	PORT(Start_ID_Cntrl : IN STD_LOGIC;
		 Update_Apk_ID : IN STD_LOGIC;
		 Reset : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 DB_K3_INP : IN STD_LOGIC;
		 DB_K2_INP : IN STD_LOGIC;
		 DB_GR1_APK_ID : IN STD_LOGIC;
		 DB_K1_INP : IN STD_LOGIC;
		 DB_K0_INP : IN STD_LOGIC;
		 DB_GR0_APK_ID : IN STD_LOGIC;
		 A_K0_D : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 A_K1_D : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 A_K2_D : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 A_K3_D : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 K1_K0_Skal : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 K3_K2_Skal : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 ID_Cntrl_Done : OUT STD_LOGIC;
		 APK_ST_ID_OK : OUT STD_LOGIC;
		 La_Ena_Skal_In : OUT STD_LOGIC;
		 La_Ena_Port_In : OUT STD_LOGIC;
		 A_nK3_ID_En : OUT STD_LOGIC;
		 A_nK2_ID_En : OUT STD_LOGIC;
		 A_nGR1_ID_Sel : OUT STD_LOGIC;
		 A_nK1_ID_En : OUT STD_LOGIC;
		 A_nK0_ID_En : OUT STD_LOGIC;
		 A_nGR0_ID_Sel : OUT STD_LOGIC;
		 K0_ID : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 K1_ID : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 K2_ID : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 K3_ID : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT chopper_pll
	PORT(inclk0 : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 c1 : OUT STD_LOGIC;
		 locked : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT skal_test
GENERIC (Gr0_16Bit : INTEGER;
			Gr0_APK_ID : INTEGER;
			Gr1_16Bit : INTEGER;
			Gr1_APK_ID : INTEGER;
			K0_Input : INTEGER;
			K0C_Def_Level : INTEGER;
			K0D_Def_Level : INTEGER;
			K1_Input : INTEGER;
			K1C_Def_Level : INTEGER;
			K1D_Def_Level : INTEGER;
			K2_Input : INTEGER;
			K2C_Def_Level : INTEGER;
			K2D_Def_Level : INTEGER;
			K3_Input : INTEGER;
			K3C_Def_Level : INTEGER;
			K3D_Def_Level : INTEGER;
			Logic_Nr_End : INTEGER;
			Logic_Nr_Start : INTEGER;
			No_Level_Test : INTEGER;
			No_Logic_Test : INTEGER;
			No_Port_Dir_Test : INTEGER;
			ST_160_Pol : INTEGER
			);
	PORT(A_K3D_SPG : IN STD_LOGIC;
		 A_K3C_SPG : IN STD_LOGIC;
		 A_K2D_SPG : IN STD_LOGIC;
		 A_K2C_SPG : IN STD_LOGIC;
		 A_K1D_SPG : IN STD_LOGIC;
		 A_K1C_SPG : IN STD_LOGIC;
		 A_K0D_SPG : IN STD_LOGIC;
		 A_K0C_SPG : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 Logik : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 St_160_Skal : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VG_Mod_Skal : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 All_Okay : OUT STD_LOGIC;
		 Mod_Skal_Ok : OUT STD_LOGIC;
		 Level_Ok : OUT STD_LOGIC;
		 Logic_Nr_Ok : OUT STD_LOGIC;
		 nK0_Switch_Ena : OUT STD_LOGIC;
		 nK1_Switch_Ena : OUT STD_LOGIC;
		 nK2_Switch_Ena : OUT STD_LOGIC;
		 nK3_Switch_Ena : OUT STD_LOGIC;
		 nSkal_Okay_Led : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT chopper_macro1
GENERIC (Clk_in_HZ : INTEGER;
			Test : INTEGER
			);
	PORT(RD_Activ : IN STD_LOGIC;
		 WR_Activ : IN STD_LOGIC;
		 Skal_OK : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 Reset : IN STD_LOGIC;
		 Off_Anforderung_In : IN STD_LOGIC;
		 Off_UU_In : IN STD_LOGIC;
		 Beam_Control_In : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Data_WR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Strahlalarm_In : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Sub_Adr_Sync : IN STD_LOGIC_VECTOR(7 DOWNTO 1);
		 Chop_m1_Rd_Activ : OUT STD_LOGIC;
		 Chop1_Macro1_Activ : OUT STD_LOGIC;
		 Chop_DT_to_MB : OUT STD_LOGIC;
		 Chop_m1_Test_Vers_Aktiv : OUT STD_LOGIC;
		 Strahlweg_Reg_WR : OUT STD_LOGIC;
		 Strahlweg_Reg_RD : OUT STD_LOGIC;
		 Strahlweg_Maske_RD : OUT STD_LOGIC;
		 Interlock_to_SE_RD : OUT STD_LOGIC;
		 Global_Status_RD : OUT STD_LOGIC;
		 Beam_Control_Out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Chop_m1_LEDs : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Chop_m1_RD_data : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Trafo_Timing_Out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT aux_signals
	PORT(beam_control_in : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 beam_control_out : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 aux_out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT kicker_leds
GENERIC (Use_LPM : INTEGER
			);
	PORT(clk : IN STD_LOGIC;
		 Led_Ena : IN STD_LOGIC;
		 Led_Sig : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 nLed_Out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT independent_clk
	PORT(		 nMaster_Clk_Ena : OUT STD_LOGIC;
		 nSlave_Clk_Ena : OUT STD_LOGIC;
		 nIndenpend_Clk_Ena : OUT STD_LOGIC;
		 Extern_Clk_OK : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT rd_apk_id
GENERIC (ST_160_Pol : INTEGER
			);
	PORT(ID_Cntrl_Done : IN STD_LOGIC;
		 Extern_Rd_Activ : IN STD_LOGIC;
		 Extern_Wr_Activ : IN STD_LOGIC;
		 Powerup_Res : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 K0_ID : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 K1_ID : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 K2_ID : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 K3_ID : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Sub_Adr_La : IN STD_LOGIC_VECTOR(7 DOWNTO 1);
		 Update_Apk_ID : OUT STD_LOGIC;
		 Rd_Apk_ID_Activ : OUT STD_LOGIC;
		 Dtack_Apk_ID : OUT STD_LOGIC;
		 Rd_Apk_ID_Port : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT rd_mux
	PORT(Sel_Chop_Out : IN STD_LOGIC;
		 Sel_Apk_ID : IN STD_LOGIC;
		 Rd_Apk_ID_Port : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Rd_Chop_Out : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Data_Rd : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT epld_vers
GENERIC (Test : INTEGER
			);
	PORT(		 Test_Activ : OUT STD_LOGIC;
		 Vers_Rev : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT kanal
	PORT(nPort_Wr : IN STD_LOGIC;
		 ID_OK : IN STD_LOGIC;
		 ID_Cntrl_Done : IN STD_LOGIC;
		 Wr_Strobe : IN STD_LOGIC;
		 Port_In_La : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 nP_CTRL : INOUT STD_LOGIC_VECTOR(2 DOWNTO 1);
		 Port_IO : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 TO_Port : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Rd_Strobe : OUT STD_LOGIC;
		 From_Port : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT k12_k23_logik_leds
GENERIC (Test : INTEGER
			);
	PORT(Logik_Aktiv : IN STD_LOGIC;
		 Test_Vers_Aktiv : IN STD_LOGIC;
		 Live_LED_In0 : IN STD_LOGIC;
		 Live_LED_In1 : IN STD_LOGIC;
		 Live_LED_In2 : IN STD_LOGIC;
		 Live_LED_In3 : IN STD_LOGIC;
		 Live_LED_In4 : IN STD_LOGIC;
		 Live_LED_In5 : IN STD_LOGIC;
		 Live_LED_In6 : IN STD_LOGIC;
		 Live_LED_In7 : IN STD_LOGIC;
		 Ena : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 Logik : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 Sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 St_160_Skal : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VG_Mod_Skal : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 nLED_Skal : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT master
	PORT(inclk0 : IN STD_LOGIC;
		 pfdena : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 c1 : OUT STD_LOGIC;
		 locked : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT modulbus_loader
GENERIC (CLK_in_Hz : INTEGER;
			I2C_Freq_in_Hz : INTEGER;
			Loader_Clk_in_Hz : INTEGER;
			LPM_Ein_ist_1 : INTEGER;
			Mod_Id : INTEGER;
			nDS_Deb_in_ns : INTEGER;
			Res_Deb_in_ns : INTEGER;
			St_160_pol : INTEGER;
			Test_Ein_ist_1 : INTEGER
			);
	PORT(Stat_IN7 : IN STD_LOGIC;
		 Stat_IN6 : IN STD_LOGIC;
		 Stat_IN5 : IN STD_LOGIC;
		 Stat_IN4 : IN STD_LOGIC;
		 Stat_IN3 : IN STD_LOGIC;
		 Stat_IN2 : IN STD_LOGIC;
		 Macro_Activ : IN STD_LOGIC;
		 Macro_Skal_Ok : IN STD_LOGIC;
		 RDnWR : IN STD_LOGIC;
		 nDS : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 nMB_Reset : IN STD_LOGIC;
		 Extern_Dtack : IN STD_LOGIC;
		 CTRL_Load : IN STD_LOGIC;
		 CTRL_Res : IN STD_LOGIC;
		 Loader_Clk : IN STD_LOGIC;
		 Loader_DB : INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Mod_Adr : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 Mod_Data : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 St_160_Auxi : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 St_160_Skal : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Sub_Adr : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 V_Data_Rd : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Vers_Rev : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VG_Mod_Adr : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 VG_Mod_Id : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VG_Mod_Skal : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 nExt_Data_En : OUT STD_LOGIC;
		 nDt_Mod_Bus : OUT STD_LOGIC;
		 Extern_Wr_Activ : OUT STD_LOGIC;
		 Extern_Wr_Fin : OUT STD_LOGIC;
		 Extern_Rd_Activ : OUT STD_LOGIC;
		 Extern_Rd_Fin : OUT STD_LOGIC;
		 Powerup_Res : OUT STD_LOGIC;
		 nInterlock : OUT STD_LOGIC;
		 ID_OK : OUT STD_LOGIC;
		 nID_OK_Led : OUT STD_LOGIC;
		 Led_Ena : OUT STD_LOGIC;
		 nPowerup_Led : OUT STD_LOGIC;
		 nDt_Led : OUT STD_LOGIC;
		 nSEL_I2C : OUT STD_LOGIC;
		 Loader_WRnRD : OUT STD_LOGIC;
		 RELOAD : OUT STD_LOGIC;
		 LOAD_OK : OUT STD_LOGIC;
		 LOAD_ERROR : OUT STD_LOGIC;
		 INIT_DONE : OUT STD_LOGIC;
		 Data_Wr_La : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Sub_Adr_La : OUT STD_LOGIC_VECTOR(7 DOWNTO 1)
	);
END COMPONENT;

SIGNAL	A_Master_Clk_Out_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	APK_Skal_Ok :  STD_LOGIC;
SIGNAL	APK_ST_ID_OK :  STD_LOGIC;
SIGNAL	Beam_Control_In :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	Beam_Control_Out :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	Chop_Dtack :  STD_LOGIC;
SIGNAL	Chop_m1_LEDs :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	Chop_m1_Rd_Activ :  STD_LOGIC;
SIGNAL	CLK :  STD_LOGIC;
SIGNAL	Data_Wr_La :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	DB_160_Skal :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DB_GR0_APK_ID :  STD_LOGIC;
SIGNAL	DB_GR1_APK_ID :  STD_LOGIC;
SIGNAL	DB_K0_INP :  STD_LOGIC;
SIGNAL	DB_K1_INP :  STD_LOGIC;
SIGNAL	DB_K2_INP :  STD_LOGIC;
SIGNAL	DB_K3_INP :  STD_LOGIC;
SIGNAL	DB_Mod_Skal :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	Dtack_Apk_ID :  STD_LOGIC;
SIGNAL	Extern_Clk :  STD_LOGIC;
SIGNAL	Extern_Clk_OK :  STD_LOGIC;
SIGNAL	Extern_Dtack :  STD_LOGIC;
SIGNAL	Extern_Rd_Activ :  STD_LOGIC;
SIGNAL	Extern_Rd_Fin :  STD_LOGIC;
SIGNAL	Extern_Wr_Activ :  STD_LOGIC;
SIGNAL	Extern_Wr_Fin :  STD_LOGIC;
SIGNAL	F_150MHz :  STD_LOGIC;
SIGNAL	ID_Cntrl_Done :  STD_LOGIC;
SIGNAL	ID_OK :  STD_LOGIC;
SIGNAL	K0_ID :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	K1_ID :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	K1_K0_Skal :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	K2_ID :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	K3_ID :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	K3_K2_Skal :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	La_Ena_Port_In :  STD_LOGIC;
SIGNAL	La_Ena_Skal_In :  STD_LOGIC;
SIGNAL	Led_Ena :  STD_LOGIC;
SIGNAL	Level_Ok :  STD_LOGIC;
SIGNAL	Logic :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	Logic_Nr_Ok :  STD_LOGIC;
SIGNAL	Mod_Skal_Ok :  STD_LOGIC;
SIGNAL	nDT_MOD_BUS :  STD_LOGIC;
SIGNAL	nInterlock :  STD_LOGIC;
SIGNAL	Powerup_Res :  STD_LOGIC;
SIGNAL	Rd_Apk_ID_Activ :  STD_LOGIC;
SIGNAL	Rd_Apk_ID_Port :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	Rd_Chop_Out :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	Skal_Okay :  STD_LOGIC;
SIGNAL	Start_ID_Cntrl :  STD_LOGIC;
SIGNAL	Strahlalarm_In :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	Sub_Adr_La :  STD_LOGIC_VECTOR(7 DOWNTO 1);
SIGNAL	Test_Activ :  STD_LOGIC;
SIGNAL	Trafo_Timing_Out :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	Update_Apk_ID :  STD_LOGIC;
SIGNAL	V_Data_Rd :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	Vers_Rev :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(0 TO 11);
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(0 TO 1);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC_VECTOR(0 TO 11);
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(0 TO 15);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(0 TO 15);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(0 TO 15);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;


BEGIN 
A_nMANUAL_RES <= '1';
RDnWR_Transceiver <= A_RDnWR;
A_nDTACKA <= SYNTHESIZED_WIRE_38;
A_nDTACKB <= SYNTHESIZED_WIRE_38;
A_nINTERLOCKA <= SYNTHESIZED_WIRE_39;
A_nINTERLOCKB <= SYNTHESIZED_WIRE_39;
A_nSRQA <= SYNTHESIZED_WIRE_40;
A_nSRQB <= SYNTHESIZED_WIRE_40;
A_nDRQB <= SYNTHESIZED_WIRE_41;
A_nDRQA <= SYNTHESIZED_WIRE_41;
SYNTHESIZED_WIRE_42 <= '0';
SYNTHESIZED_WIRE_43 <= "000000000000";
SYNTHESIZED_WIRE_44 <= '0';
SYNTHESIZED_WIRE_45 <= '0';
SYNTHESIZED_WIRE_46 <= "00";
SYNTHESIZED_WIRE_47 <= '0';
SYNTHESIZED_WIRE_48 <= "000000000000";
SYNTHESIZED_WIRE_25 <= "1111111111111111";
SYNTHESIZED_WIRE_26 <= '1';
SYNTHESIZED_WIRE_27 <= "0000000000000000";
SYNTHESIZED_WIRE_28 <= '1';
SYNTHESIZED_WIRE_29 <= "0000000000000000";
SYNTHESIZED_WIRE_30 <= '1';
SYNTHESIZED_WIRE_31 <= '1';
SYNTHESIZED_WIRE_49 <= '0';
SYNTHESIZED_WIRE_34 <= '1';
SYNTHESIZED_WIRE_50 <= '0';



b2v_Bus_IO_inst : bus_io
GENERIC MAP(I0_1_is_Input => 1,
			I0_2_is_Input => 1,
			I0_3_is_Input => 1,
			I0_4_is_Input => 1,
			I0_5_is_Input => 1,
			ST_160_Pol => 1
			)
PORT MAP(To_IO_5 => SYNTHESIZED_WIRE_42,
		 To_IO_4 => SYNTHESIZED_WIRE_42,
		 To_IO_3 => SYNTHESIZED_WIRE_42,
		 To_IO_2 => SYNTHESIZED_WIRE_42,
		 To_IO_1 => SYNTHESIZED_WIRE_42,
		 A_Bus_IO => A_Bus_IO);


b2v_DB_Skal : debounce_skal
GENERIC MAP(Clk_in_Hz => 20000000,
			DB_in_ns => 200,
			Test => 0
			)
PORT MAP(A_VG_K1_INP => A_VG_K1_INP,
		 A_VG_K0_INP => A_VG_K0_INP,
		 A_GR0_APK_ID => A_GR0_APK_ID,
		 A_GR0_16BIT => A_GR0_16BIT,
		 A_VG_K3_INP => A_VG_K3_INP,
		 A_VG_K2_INP => A_VG_K2_INP,
		 A_GR1_APK_ID => A_GR1_APK_ID,
		 A_GR1_16BIT => A_GR1_16BIT,
		 Latch_Inputs => La_Ena_Skal_In,
		 Reset => Powerup_Res,
		 clk => A_Master_Clk_Out_ALTERA_SYNTHESIZED,
		 A_VG_K0_MOD => A_VG_K0_MOD,
		 A_VG_K1_MOD => A_VG_K1_MOD,
		 A_VG_K2_MOD => A_VG_K2_MOD,
		 A_VG_K3_MOD => A_VG_K3_MOD,
		 Logic => A_VG_Log_ID,
		 DB_K1_INP => DB_K1_INP,
		 DB_K0_INP => DB_K0_INP,
		 DB_GR0_APK_ID => DB_GR0_APK_ID,
		 DB_K3_INP => DB_K3_INP,
		 DB_K2_INP => DB_K2_INP,
		 DB_GR1_APK_ID => DB_GR1_APK_ID,
		 DB_Valid => Start_ID_Cntrl,
		 DB_160_Skal => DB_160_Skal,
		 DB_Logic => Logic,
		 DB_Mod_Skal => DB_Mod_Skal,
		 K1_K0_Skal => K1_K0_Skal,
		 K3_K2_Skal => K3_K2_Skal);


b2v_ID_Cntrl : apk_stecker_id_cntrl
GENERIC MAP(Clk_in_Hz => 150000000,
			K0_APK_ST_ID => 53312,
			K1_APK_ST_ID => 53319,
			K2_APK_ST_ID => 60720,
			K3_APK_ST_ID => 60720,
			ST_160_Pol => 1,
			Use_LPM => 1,
			Wait_in_ns => 200
			)
PORT MAP(Start_ID_Cntrl => Start_ID_Cntrl,
		 Update_Apk_ID => Update_Apk_ID,
		 Reset => Powerup_Res,
		 clk => F_150MHz,
		 DB_K3_INP => DB_K3_INP,
		 DB_K2_INP => DB_K2_INP,
		 DB_GR1_APK_ID => DB_GR1_APK_ID,
		 DB_K1_INP => DB_K1_INP,
		 DB_K0_INP => DB_K0_INP,
		 DB_GR0_APK_ID => DB_GR0_APK_ID,
		 A_K0_D => A_K0_D,
		 A_K1_D => A_K1_D,
		 A_K2_D => A_K2_D,
		 A_K3_D => A_K3_D,
		 K1_K0_Skal => K1_K0_Skal,
		 K3_K2_Skal => K3_K2_Skal,
		 ID_Cntrl_Done => ID_Cntrl_Done,
		 APK_ST_ID_OK => APK_ST_ID_OK,
		 La_Ena_Skal_In => La_Ena_Skal_In,
		 La_Ena_Port_In => La_Ena_Port_In,
		 A_nK3_ID_En => A_nK3_ID_EN,
		 A_nK2_ID_En => A_nK2_ID_EN,
		 A_nGR1_ID_Sel => A_nGR1_ID_SEL,
		 A_nK1_ID_En => A_nK1_ID_EN,
		 A_nK0_ID_En => A_nK0_ID_EN,
		 A_nGR0_ID_Sel => A_nGR0_ID_SEL,
		 K0_ID => K0_ID,
		 K1_ID => K1_ID,
		 K2_ID => K2_ID,
		 K3_ID => K3_ID);


APK_Skal_Ok <= Skal_Okay AND APK_ST_ID_OK;


b2v_inst1 : chopper_pll
PORT MAP(inclk0 => Chopper_Clk,
		 c0 => CLK);



PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(0) = '1') THEN
	TP(12) <= SYNTHESIZED_WIRE_43(0);
ELSE
	TP(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(1) = '1') THEN
	TP(11) <= SYNTHESIZED_WIRE_43(1);
ELSE
	TP(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(2) = '1') THEN
	TP(10) <= SYNTHESIZED_WIRE_43(2);
ELSE
	TP(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(3) = '1') THEN
	TP(9) <= SYNTHESIZED_WIRE_43(3);
ELSE
	TP(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(4) = '1') THEN
	TP(8) <= SYNTHESIZED_WIRE_43(4);
ELSE
	TP(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(5) = '1') THEN
	TP(7) <= SYNTHESIZED_WIRE_43(5);
ELSE
	TP(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(6) = '1') THEN
	TP(6) <= SYNTHESIZED_WIRE_43(6);
ELSE
	TP(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(7) = '1') THEN
	TP(5) <= SYNTHESIZED_WIRE_43(7);
ELSE
	TP(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(8) = '1') THEN
	TP(4) <= SYNTHESIZED_WIRE_43(8);
ELSE
	TP(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(9) = '1') THEN
	TP(3) <= SYNTHESIZED_WIRE_43(9);
ELSE
	TP(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(10) = '1') THEN
	TP(2) <= SYNTHESIZED_WIRE_43(10);
ELSE
	TP(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_43,SYNTHESIZED_WIRE_43)
BEGIN
if (SYNTHESIZED_WIRE_43(11) = '1') THEN
	TP(1) <= SYNTHESIZED_WIRE_43(11);
ELSE
	TP(1) <= 'Z';
END IF;
END PROCESS;



b2v_inst11 : skal_test
GENERIC MAP(Gr0_16Bit => 1,
			Gr0_APK_ID => 1,
			Gr1_16Bit => 1,
			Gr1_APK_ID => 1,
			K0_Input => 1,
			K0C_Def_Level => 1,
			K0D_Def_Level => 0,
			K1_Input => 1,
			K1C_Def_Level => 1,
			K1D_Def_Level => 0,
			K2_Input => 0,
			K2C_Def_Level => 1,
			K2D_Def_Level => 0,
			K3_Input => 0,
			K3C_Def_Level => 1,
			K3D_Def_Level => 0,
			Logic_Nr_End => 1,
			Logic_Nr_Start => 1,
			No_Level_Test => 0,
			No_Logic_Test => 0,
			No_Port_Dir_Test => 0,
			ST_160_Pol => 1
			)
PORT MAP(A_K3D_SPG => A_K3D_SPG,
		 A_K3C_SPG => A_K3C_SPG,
		 A_K2D_SPG => A_K2D_SPG,
		 A_K2C_SPG => A_K2C_SPG,
		 A_K1D_SPG => A_K1D_SPG,
		 A_K1C_SPG => A_K1C_SPG,
		 A_K0D_SPG => A_K0D_SPG,
		 A_K0C_SPG => A_K0C_SPG,
		 clk => CLK,
		 Logik => Logic,
		 St_160_Skal => DB_160_Skal,
		 VG_Mod_Skal => DB_Mod_Skal,
		 All_Okay => Skal_Okay,
		 Mod_Skal_Ok => Mod_Skal_Ok,
		 Level_Ok => Level_Ok,
		 Logic_Nr_Ok => Logic_Nr_Ok,
		 nK0_Switch_Ena => nK0_SWITCH_ENA,
		 nK1_Switch_Ena => nK1_SWITCH_ENA,
		 nK2_Switch_Ena => nK2_SWITCH_ENA,
		 nK3_Switch_Ena => nK3_SWITCH_ENA,
		 nSkal_Okay_Led => nSkal_OK_Led);


PROCESS(SYNTHESIZED_WIRE_44,SYNTHESIZED_WIRE_44)
BEGIN
if (SYNTHESIZED_WIRE_44 = '1') THEN
	A_AUX_CA <= SYNTHESIZED_WIRE_44;
ELSE
	A_AUX_CA <= 'Z';
END IF;
END PROCESS;



PROCESS(SYNTHESIZED_WIRE_45,SYNTHESIZED_WIRE_45)
BEGIN
if (SYNTHESIZED_WIRE_45 = '1') THEN
	A_AUX_CB <= SYNTHESIZED_WIRE_45;
ELSE
	A_AUX_CB <= 'Z';
END IF;
END PROCESS;



b2v_inst12 : chopper_macro1
GENERIC MAP(Clk_in_HZ => 200000000,
			Test => 0
			)
PORT MAP(RD_Activ => Extern_Rd_Activ,
		 WR_Activ => Extern_Wr_Activ,
		 Skal_OK => APK_Skal_Ok,
		 Clk => CLK,
		 Reset => Powerup_Res,
		 Off_Anforderung_In => A_Bus_IO(1),
		 Off_UU_In => A_Bus_IO(2),
		 Beam_Control_In => Beam_Control_In,
		 Data_WR => Data_Wr_La,
		 Strahlalarm_In => Strahlalarm_In,
		 Sub_Adr_Sync => Sub_Adr_La,
		 Chop_m1_Rd_Activ => Chop_m1_Rd_Activ,
		 Chop_DT_to_MB => Chop_Dtack,
		 Beam_Control_Out => Beam_Control_Out,
		 Chop_m1_LEDs => Chop_m1_LEDs,
		 Chop_m1_RD_data => Rd_Chop_Out,
		 Trafo_Timing_Out => Trafo_Timing_Out);


b2v_inst13 : aux_signals
PORT MAP(beam_control_in => Beam_Control_In,
		 beam_control_out => Beam_Control_Out,
		 aux_out => SYNTHESIZED_WIRE_24);



b2v_inst17 : kicker_leds
GENERIC MAP(Use_LPM => 1
			)
PORT MAP(clk => CLK,
		 Led_Ena => Led_Ena,
		 Led_Sig => Chop_m1_LEDs,
		 nLed_Out => nLED);

SYNTHESIZED_WIRE_38 <= nDT_MOD_BUS;



b2v_inst2 : independent_clk
PORT MAP(		 nMaster_Clk_Ena => nMaster_Clk_ENA,
		 nSlave_Clk_Ena => nSlave_Clk_ENA,
		 nIndenpend_Clk_Ena => nIndepend_Clk_Ena,
		 Extern_Clk_OK => Extern_Clk_OK);










SYNTHESIZED_WIRE_12 <= NOT(SYNTHESIZED_WIRE_46);



b2v_inst4 : rd_apk_id
GENERIC MAP(ST_160_Pol => 1
			)
PORT MAP(ID_Cntrl_Done => ID_Cntrl_Done,
		 Extern_Rd_Activ => Extern_Rd_Activ,
		 Extern_Wr_Activ => Extern_Wr_Activ,
		 Powerup_Res => Powerup_Res,
		 Clk => CLK,
		 K0_ID => K0_ID,
		 K1_ID => K1_ID,
		 K2_ID => K2_ID,
		 K3_ID => K3_ID,
		 Sub_Adr_La => Sub_Adr_La,
		 Update_Apk_ID => Update_Apk_ID,
		 Rd_Apk_ID_Activ => Rd_Apk_ID_Activ,
		 Dtack_Apk_ID => Dtack_Apk_ID,
		 Rd_Apk_ID_Port => Rd_Apk_ID_Port);



Extern_Dtack <= Dtack_Apk_ID OR Chop_Dtack;



b2v_inst6 : rd_mux
PORT MAP(Sel_Chop_Out => Chop_m1_Rd_Activ,
		 Sel_Apk_ID => Rd_Apk_ID_Activ,
		 Rd_Apk_ID_Port => Rd_Apk_ID_Port,
		 Rd_Chop_Out => Rd_Chop_Out,
		 Data_Rd => V_Data_Rd);


PROCESS(SYNTHESIZED_WIRE_12,SYNTHESIZED_WIRE_46)
BEGIN
if (SYNTHESIZED_WIRE_46(0) = '1') THEN
	A_VG_IO_Res(1) <= SYNTHESIZED_WIRE_12(1);
ELSE
	A_VG_IO_Res(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_12,SYNTHESIZED_WIRE_46)
BEGIN
if (SYNTHESIZED_WIRE_46(1) = '1') THEN
	A_VG_IO_Res(0) <= SYNTHESIZED_WIRE_12(0);
ELSE
	A_VG_IO_Res(0) <= 'Z';
END IF;
END PROCESS;


b2v_inst7 : epld_vers
GENERIC MAP(Test => 0
			)
PORT MAP(		 Test_Activ => Test_Activ,
		 Vers_Rev => Vers_Rev);



PROCESS(SYNTHESIZED_WIRE_47,SYNTHESIZED_WIRE_47)
BEGIN
if (SYNTHESIZED_WIRE_47 = '1') THEN
	SYNTHESIZED_WIRE_40 <= SYNTHESIZED_WIRE_47;
ELSE
	SYNTHESIZED_WIRE_40 <= 'Z';
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_47,SYNTHESIZED_WIRE_47)
BEGIN
if (SYNTHESIZED_WIRE_47 = '1') THEN
	SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_47;
ELSE
	SYNTHESIZED_WIRE_41 <= 'Z';
END IF;
END PROCESS;

SYNTHESIZED_WIRE_39 <= nInterlock;



PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(0) = '1') THEN
	A_AUX_A(11) <= SYNTHESIZED_WIRE_48(0);
ELSE
	A_AUX_A(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(1) = '1') THEN
	A_AUX_A(10) <= SYNTHESIZED_WIRE_48(1);
ELSE
	A_AUX_A(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(2) = '1') THEN
	A_AUX_A(9) <= SYNTHESIZED_WIRE_48(2);
ELSE
	A_AUX_A(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(3) = '1') THEN
	A_AUX_A(8) <= SYNTHESIZED_WIRE_48(3);
ELSE
	A_AUX_A(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(4) = '1') THEN
	A_AUX_A(7) <= SYNTHESIZED_WIRE_48(4);
ELSE
	A_AUX_A(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(5) = '1') THEN
	A_AUX_A(6) <= SYNTHESIZED_WIRE_48(5);
ELSE
	A_AUX_A(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(6) = '1') THEN
	A_AUX_A(5) <= SYNTHESIZED_WIRE_48(6);
ELSE
	A_AUX_A(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(7) = '1') THEN
	A_AUX_A(4) <= SYNTHESIZED_WIRE_48(7);
ELSE
	A_AUX_A(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(8) = '1') THEN
	A_AUX_A(3) <= SYNTHESIZED_WIRE_48(8);
ELSE
	A_AUX_A(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(9) = '1') THEN
	A_AUX_A(2) <= SYNTHESIZED_WIRE_48(9);
ELSE
	A_AUX_A(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(10) = '1') THEN
	A_AUX_A(1) <= SYNTHESIZED_WIRE_48(10);
ELSE
	A_AUX_A(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(11) = '1') THEN
	A_AUX_A(0) <= SYNTHESIZED_WIRE_48(11);
ELSE
	A_AUX_A(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(0) = '1') THEN
	A_AUX_B(11) <= SYNTHESIZED_WIRE_48(0);
ELSE
	A_AUX_B(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(1) = '1') THEN
	A_AUX_B(10) <= SYNTHESIZED_WIRE_48(1);
ELSE
	A_AUX_B(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(2) = '1') THEN
	A_AUX_B(9) <= SYNTHESIZED_WIRE_48(2);
ELSE
	A_AUX_B(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(3) = '1') THEN
	A_AUX_B(8) <= SYNTHESIZED_WIRE_48(3);
ELSE
	A_AUX_B(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(4) = '1') THEN
	A_AUX_B(7) <= SYNTHESIZED_WIRE_48(4);
ELSE
	A_AUX_B(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(5) = '1') THEN
	A_AUX_B(6) <= SYNTHESIZED_WIRE_48(5);
ELSE
	A_AUX_B(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(6) = '1') THEN
	A_AUX_B(5) <= SYNTHESIZED_WIRE_48(6);
ELSE
	A_AUX_B(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(7) = '1') THEN
	A_AUX_B(4) <= SYNTHESIZED_WIRE_48(7);
ELSE
	A_AUX_B(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(8) = '1') THEN
	A_AUX_B(3) <= SYNTHESIZED_WIRE_48(8);
ELSE
	A_AUX_B(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(9) = '1') THEN
	A_AUX_B(2) <= SYNTHESIZED_WIRE_48(9);
ELSE
	A_AUX_B(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(10) = '1') THEN
	A_AUX_B(1) <= SYNTHESIZED_WIRE_48(10);
ELSE
	A_AUX_B(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(11) = '1') THEN
	A_AUX_B(0) <= SYNTHESIZED_WIRE_48(11);
ELSE
	A_AUX_B(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(0) = '1') THEN
	A_AUX_C(11) <= SYNTHESIZED_WIRE_48(0);
ELSE
	A_AUX_C(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(1) = '1') THEN
	A_AUX_C(10) <= SYNTHESIZED_WIRE_48(1);
ELSE
	A_AUX_C(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(2) = '1') THEN
	A_AUX_C(9) <= SYNTHESIZED_WIRE_48(2);
ELSE
	A_AUX_C(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(3) = '1') THEN
	A_AUX_C(8) <= SYNTHESIZED_WIRE_48(3);
ELSE
	A_AUX_C(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(4) = '1') THEN
	A_AUX_C(7) <= SYNTHESIZED_WIRE_48(4);
ELSE
	A_AUX_C(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(5) = '1') THEN
	A_AUX_C(6) <= SYNTHESIZED_WIRE_48(5);
ELSE
	A_AUX_C(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(6) = '1') THEN
	A_AUX_C(5) <= SYNTHESIZED_WIRE_48(6);
ELSE
	A_AUX_C(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(7) = '1') THEN
	A_AUX_C(4) <= SYNTHESIZED_WIRE_48(7);
ELSE
	A_AUX_C(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(8) = '1') THEN
	A_AUX_C(3) <= SYNTHESIZED_WIRE_48(8);
ELSE
	A_AUX_C(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(9) = '1') THEN
	A_AUX_C(2) <= SYNTHESIZED_WIRE_48(9);
ELSE
	A_AUX_C(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(10) = '1') THEN
	A_AUX_C(1) <= SYNTHESIZED_WIRE_48(10);
ELSE
	A_AUX_C(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_48)
BEGIN
if (SYNTHESIZED_WIRE_48(11) = '1') THEN
	A_AUX_C(0) <= SYNTHESIZED_WIRE_48(11);
ELSE
	A_AUX_C(0) <= 'Z';
END IF;
END PROCESS;




PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(0) = '1') THEN
	A_Test(15) <= SYNTHESIZED_WIRE_24(15);
ELSE
	A_Test(15) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(1) = '1') THEN
	A_Test(14) <= SYNTHESIZED_WIRE_24(14);
ELSE
	A_Test(14) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(2) = '1') THEN
	A_Test(13) <= SYNTHESIZED_WIRE_24(13);
ELSE
	A_Test(13) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(3) = '1') THEN
	A_Test(12) <= SYNTHESIZED_WIRE_24(12);
ELSE
	A_Test(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(4) = '1') THEN
	A_Test(11) <= SYNTHESIZED_WIRE_24(11);
ELSE
	A_Test(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(5) = '1') THEN
	A_Test(10) <= SYNTHESIZED_WIRE_24(10);
ELSE
	A_Test(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(6) = '1') THEN
	A_Test(9) <= SYNTHESIZED_WIRE_24(9);
ELSE
	A_Test(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(7) = '1') THEN
	A_Test(8) <= SYNTHESIZED_WIRE_24(8);
ELSE
	A_Test(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(8) = '1') THEN
	A_Test(7) <= SYNTHESIZED_WIRE_24(7);
ELSE
	A_Test(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(9) = '1') THEN
	A_Test(6) <= SYNTHESIZED_WIRE_24(6);
ELSE
	A_Test(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(10) = '1') THEN
	A_Test(5) <= SYNTHESIZED_WIRE_24(5);
ELSE
	A_Test(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(11) = '1') THEN
	A_Test(4) <= SYNTHESIZED_WIRE_24(4);
ELSE
	A_Test(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(12) = '1') THEN
	A_Test(3) <= SYNTHESIZED_WIRE_24(3);
ELSE
	A_Test(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(13) = '1') THEN
	A_Test(2) <= SYNTHESIZED_WIRE_24(2);
ELSE
	A_Test(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(14) = '1') THEN
	A_Test(1) <= SYNTHESIZED_WIRE_24(1);
ELSE
	A_Test(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
if (SYNTHESIZED_WIRE_25(15) = '1') THEN
	A_Test(0) <= SYNTHESIZED_WIRE_24(0);
ELSE
	A_Test(0) <= 'Z';
END IF;
END PROCESS;


b2v_K0 : kanal
PORT MAP(nPort_Wr => DB_K0_INP,
		 ID_OK => ID_OK,
		 ID_Cntrl_Done => ID_Cntrl_Done,
		 Wr_Strobe => SYNTHESIZED_WIRE_26,
		 Port_In_La => La_Ena_Port_In,
		 clk => CLK,
		 nP_CTRL => A_nK0_CTRL,
		 Port_IO => A_K0_D,
		 TO_Port => SYNTHESIZED_WIRE_27,
		 From_Port => Beam_Control_In);


b2v_K1 : kanal
PORT MAP(nPort_Wr => DB_K1_INP,
		 ID_OK => ID_OK,
		 ID_Cntrl_Done => ID_Cntrl_Done,
		 Wr_Strobe => SYNTHESIZED_WIRE_28,
		 Port_In_La => La_Ena_Port_In,
		 clk => CLK,
		 nP_CTRL => A_nK1_CTRL,
		 Port_IO => A_K1_D,
		 TO_Port => SYNTHESIZED_WIRE_29,
		 From_Port => Strahlalarm_In);


b2v_K2 : kanal
PORT MAP(nPort_Wr => DB_K2_INP,
		 ID_OK => ID_OK,
		 ID_Cntrl_Done => ID_Cntrl_Done,
		 Wr_Strobe => SYNTHESIZED_WIRE_30,
		 Port_In_La => La_Ena_Port_In,
		 clk => CLK,
		 nP_CTRL => A_nK2_CTRL,
		 Port_IO => A_K2_D,
		 TO_Port => Trafo_Timing_Out);


b2v_K3 : kanal
PORT MAP(nPort_Wr => DB_K3_INP,
		 ID_OK => ID_OK,
		 ID_Cntrl_Done => ID_Cntrl_Done,
		 Wr_Strobe => SYNTHESIZED_WIRE_31,
		 Port_In_La => La_Ena_Port_In,
		 clk => CLK,
		 nP_CTRL => A_nK3_CTRL,
		 Port_IO => A_K3_D,
		 TO_Port => Beam_Control_Out);


b2v_Logik_Leds : k12_k23_logik_leds
GENERIC MAP(Test => 0
			)
PORT MAP(Logik_Aktiv => Skal_Okay,
		 Test_Vers_Aktiv => Test_Activ,
		 Live_LED_In0 => Extern_Clk_OK,
		 Live_LED_In1 => SYNTHESIZED_WIRE_49,
		 Live_LED_In2 => SYNTHESIZED_WIRE_49,
		 Live_LED_In3 => APK_ST_ID_OK,
		 Live_LED_In4 => Logic_Nr_Ok,
		 Live_LED_In5 => Level_Ok,
		 Live_LED_In6 => Mod_Skal_Ok,
		 Live_LED_In7 => Skal_Okay,
		 Ena => Led_Ena,
		 clk => CLK,
		 Logik => Logic,
		 Sel => nSEL_LED_GRP,
		 St_160_Skal => DB_160_Skal,
		 VG_Mod_Skal => DB_Mod_Skal,
		 nLED_Skal => nLED_Skal);


b2v_master_clk1 : master
PORT MAP(inclk0 => F_TCXO_In,
		 pfdena => SYNTHESIZED_WIRE_34,
		 c0 => A_Master_Clk_Out_ALTERA_SYNTHESIZED,
		 c1 => F_150MHz);


b2v_MB_Ld : modulbus_loader
GENERIC MAP(CLK_in_Hz => 200000000,
			I2C_Freq_in_Hz => 400000,
			Loader_Clk_in_Hz => 150000000,
			LPM_Ein_ist_1 => 1,
			Mod_Id => 39,
			nDS_Deb_in_ns => 80,
			Res_Deb_in_ns => 100,
			St_160_pol => 1,
			Test_Ein_ist_1 => 0
			)
PORT MAP(Stat_IN7 => Skal_Okay,
		 Stat_IN6 => Mod_Skal_Ok,
		 Stat_IN5 => Level_Ok,
		 Stat_IN4 => Logic_Nr_Ok,
		 Stat_IN3 => APK_ST_ID_OK,
		 Stat_IN2 => SYNTHESIZED_WIRE_50,
		 Macro_Activ => SYNTHESIZED_WIRE_50,
		 Macro_Skal_Ok => SYNTHESIZED_WIRE_50,
		 RDnWR => A_RDnWR,
		 nDS => A_nDS,
		 CLK => CLK,
		 nMB_Reset => A_nMB_Reset,
		 Extern_Dtack => Extern_Dtack,
		 CTRL_Load => CTRL_LOAD,
		 CTRL_Res => CTRL_RES,
		 Loader_Clk => F_150MHz,
		 Loader_DB => Loader_DB,
		 Mod_Adr => A_A,
		 Mod_Data => A_Mod_Data,
		 St_160_Auxi => Logic,
		 St_160_Skal => DB_160_Skal,
		 Sub_Adr => A_Sub_Adr,
		 V_Data_Rd => V_Data_Rd,
		 Vers_Rev => Vers_Rev,
		 VG_Mod_Adr => A_VG_A,
		 VG_Mod_Id => A_VG_ID,
		 VG_Mod_Skal => DB_Mod_Skal,
		 nExt_Data_En => nExt_Data_En,
		 nDt_Mod_Bus => nDT_MOD_BUS,
		 Extern_Wr_Activ => Extern_Wr_Activ,
		 Extern_Rd_Activ => Extern_Rd_Activ,
		 Powerup_Res => Powerup_Res,
		 nInterlock => nInterlock,
		 ID_OK => ID_OK,
		 nID_OK_Led => nID_OK_Led,
		 Led_Ena => Led_Ena,
		 nPowerup_Led => nPowerup_Led,
		 nDt_Led => nDT_Led,
		 nSEL_I2C => A_I2C_SCL,
		 Loader_WRnRD => Loader_WRnRD,
		 RELOAD => RELOAD,
		 LOAD_OK => LOAD_OK,
		 LOAD_ERROR => LOAD_ERROR,
		 INIT_DONE => INIT_DONE,
		 Data_Wr_La => Data_Wr_La,
		 Sub_Adr_La => Sub_Adr_La);

A_Master_Clk_Out <= A_Master_Clk_Out_ALTERA_SYNTHESIZED;

END bdf_type;