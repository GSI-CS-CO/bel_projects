-- megafunction wizard: %ALTASMI_PARALLEL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTASMI_PARALLEL 

-- ============================================================
-- File Name: altasmi.vhd
-- Megafunction Name(s):
-- 			ALTASMI_PARALLEL
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Standard Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altasmi_parallel CBX_AUTO_BLACKBOX="ALL" DATA_WIDTH="STANDARD" DEVICE_FAMILY="Arria II GX" ENABLE_SIM="FALSE" EPCS_TYPE="EPCS128" FLASH_RSTPIN="FALSE" PAGE_SIZE=256 PORT_BULK_ERASE="PORT_UNUSED" PORT_DIE_ERASE="PORT_UNUSED" PORT_EN4B_ADDR="PORT_UNUSED" PORT_EX4B_ADDR="PORT_UNUSED" PORT_FAST_READ="PORT_USED" PORT_ILLEGAL_ERASE="PORT_USED" PORT_ILLEGAL_WRITE="PORT_USED" PORT_RDID_OUT="PORT_USED" PORT_READ_ADDRESS="PORT_USED" PORT_READ_DUMMYCLK="PORT_UNUSED" PORT_READ_RDID="PORT_USED" PORT_READ_SID="PORT_UNUSED" PORT_READ_STATUS="PORT_USED" PORT_SECTOR_ERASE="PORT_USED" PORT_SECTOR_PROTECT="PORT_UNUSED" PORT_SHIFT_BYTES="PORT_USED" PORT_WREN="PORT_UNUSED" PORT_WRITE="PORT_USED" USE_ASMIBLOCK="OFF" USE_EAB="ON" WRITE_DUMMY_CLK=0 addr asmi_dataoe asmi_dataout asmi_dclk asmi_scein asmi_sdoin busy clkin data_valid datain dataout fast_read illegal_erase illegal_write rden rdid_out read_address read_rdid read_status reset sector_erase shift_bytes status_out write INTENDED_DEVICE_FAMILY="Arria II GX" ALTERA_INTERNAL_OPTIONS=SUPPRESS_DA_RULE_INTERNAL=C106
--VERSION_BEGIN 18.1 cbx_a_gray2bin 2018:09:12:13:04:09:SJ cbx_a_graycounter 2018:09:12:13:04:09:SJ cbx_altasmi_parallel 2018:09:12:13:04:09:SJ cbx_altdpram 2018:09:12:13:04:09:SJ cbx_altera_counter 2018:09:12:13:04:09:SJ cbx_altera_syncram 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_arriav 2018:09:12:13:04:09:SJ cbx_cyclone 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_fifo_common 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_counter 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_nightfury 2018:09:12:13:04:09:SJ cbx_scfifo 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ cbx_zippleback 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = a_graycounter 4 lpm_compare 2 lpm_counter 3 lut 29 mux21 2 reg 152 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altasmi_altasmi_parallel_di43 IS 
	 PORT 
	 ( 
		 addr	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 asmi_dataoe	:	OUT  STD_LOGIC;
		 asmi_dataout	:	IN  STD_LOGIC := '0';
		 asmi_dclk	:	OUT  STD_LOGIC;
		 asmi_scein	:	OUT  STD_LOGIC;
		 asmi_sdoin	:	OUT  STD_LOGIC;
		 busy	:	OUT  STD_LOGIC;
		 clkin	:	IN  STD_LOGIC;
		 data_valid	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 fast_read	:	IN  STD_LOGIC := '0';
		 illegal_erase	:	OUT  STD_LOGIC;
		 illegal_write	:	OUT  STD_LOGIC;
		 rden	:	IN  STD_LOGIC;
		 rdid_out	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 read_address	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 read_rdid	:	IN  STD_LOGIC := '0';
		 read_status	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC := '0';
		 sector_erase	:	IN  STD_LOGIC := '0';
		 shift_bytes	:	IN  STD_LOGIC := '0';
		 status_out	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 write	:	IN  STD_LOGIC := '0'
	 ); 
 END altasmi_altasmi_parallel_di43;

 ARCHITECTURE RTL OF altasmi_altasmi_parallel_di43 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "SUPPRESS_DA_RULE_INTERNAL=C106";

	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range174w179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range177w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_addbyte_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_end_operation114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range126w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range124w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_end1_cyc_reg_in_wire57w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w367w368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range116w119w364w365w366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range116w119w369w370w371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range116w117w118w378w379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w121w454w455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w119w364w365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w119w389w390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w119w369w370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w117w118w378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range116w121w454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range116w119w364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range116w119w389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range116w119w369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range116w119w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range116w119w362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range115w120w138w139w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range115w120w138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range116w117w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range116w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range116w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range115w120w138w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range115w120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range116w117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w110w111w112w113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w_q_range115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_q_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_lg_w_q_range655w656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_lg_w_q_range653w654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w648w649w650w651w652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_wrstage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_q_range653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_q_range655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 add_msb_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_add_msb_reg_ena	:	STD_LOGIC;
	 SIGNAL	 add_rollover_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 addr_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range428w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_asmi_opcode_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 asmi_opcode_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_asmi_opcode_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_asmi_opcode_reg_w_q_range184w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 buf_empty_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 busy_delay_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 busy_det_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rdid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rstat_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_write_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cnt_bfend_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 do_wrmemadd_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dvalid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dvalid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_dvalid_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 dvalid_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_hdlyreg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_pgwrop_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_pgwrop_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_rbyte_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_rbyte_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_end_rbyte_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 end_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 fast_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_fast_read_reg_ena	:	STD_LOGIC;
	 SIGNAL	 ill_erase_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ill_write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 illegal_erase_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 illegal_write_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 illegal_write_prot_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_cnt_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 maxcnt_shift_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 maxcnt_shift_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ncs_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_ncs_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_ncs_reg_w_lg_q415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_pgwrbuf_dataout_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 pgwrbuf_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_pgwrbuf_dataout_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_pgwrbuf_dataout_w_q_range596w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 power_up_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rdid_out_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_add_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 read_add_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_add_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL	 read_bufdly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_data_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_read_dout_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_dout_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_dout_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 read_rdid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_rdid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 read_status_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_status_reg_ena	:	STD_LOGIC;
	 SIGNAL	 sec_erase_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_sec_erase_reg_ena	:	STD_LOGIC;
	 SIGNAL	 shftpgwr_data_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage2_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage4_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 start_wrpoll_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_start_wrpoll_reg_ena	:	STD_LOGIC;
	 SIGNAL	 start_wrpoll_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_int_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 statreg_int	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_int_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_statreg_out_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 statreg_out	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_out_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 write_prot_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_write_prot_reg_ena	:	STD_LOGIC;
	 SIGNAL	 write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_write_reg_ena	:	STD_LOGIC;
	 SIGNAL	 write_rstat_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cmpr4_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr4_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr4_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr5_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr5_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_q	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_read_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_read_buf789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_read_cntr_q	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire516w517w518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_data	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_q	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_rden_wire516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	wire_mux211_dataout	:	STD_LOGIC;
	 SIGNAL	wire_mux212_dataout	:	STD_LOGIC;
	 SIGNAL  wire_scfifo3_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_scfifo3_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_scfifo3_rdreq	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_read_buf593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_scfifo3_wrreq	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_shift_bytes_wire591w592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_scfifo3_w_q_range599w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_scfifo3_w_q_range604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w568w569w570w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w568w569w570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w814w815w816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w568w569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w814w815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w243w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w236w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_end_ophdly564w565w566w567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode200w201w202w287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode200w201w202w203w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode239w240w241w242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode210w211w212w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode210w211w212w213w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode251w252w253w309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode251w252w253w254w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode232w233w234w235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read394w395w396w397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write563w811w812w813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w661w806w807w817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read335w507w508w509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase68w450w451w452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_end_ophdly564w565w566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode200w201w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode205w206w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode215w220w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode215w220w221w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode215w216w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode215w216w217w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode239w240w241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode210w211w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode251w252w253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode232w233w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp2_wire677w678w679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp2_wire677w678w682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp2_wire677w684w685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp2_wire677w684w687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read394w395w396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read394w395w453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write563w811w812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w661w806w807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read335w507w508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_erase68w450w451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire689w690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire689w692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire694w695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire694w697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_4baddr192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_ex4baddr187w188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_polling577w578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write223w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write77w373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_ophdly564w565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_read_byte514w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode194w283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode194w195w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode189w281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode189w190w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode225w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode225w226w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode200w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode205w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode245w305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode245w246w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode248w307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode248w249w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode228w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode228w229w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode256w311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode256w257w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode259w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode259w260w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode215w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode215w216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode239w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode210w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode251w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode197w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode197w198w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode232w233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_reach_max_cnt643w644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage3_wire59w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_start_poll380w381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire677w678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire677w684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read394w395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write563w811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly597w598w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w648w649w650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w661w806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write86w87w442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read335w507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase68w450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_operation579w580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rden_wire446w447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie427w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp2_wire689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp2_wire694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_nonvolatile360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_ophdly564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read_byte514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_in_operation52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy431w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_reach_max_cnt643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly600w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_opcode185w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire429w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_start_poll380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range699w712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range702w719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range704w724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range706w729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range708w734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range710w738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write77w392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire350w351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_stage4_wire336w337w338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_stat346w347w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp0_wire675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp1_wire676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp2_wire677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_buf_empty780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_busy_wire3w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clkin_wire48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_rstat_wire50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_sid_wire49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_die_erase561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_fast_read393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_memadd459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_nonvolatile10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_volatile231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_prot559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write_volatile238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_add_cycle97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_fast_read91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_ophdly51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_pgwr_data76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reach_max_cnt607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_rdid_wire14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_sid_wire13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_status_wire29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sec_protect_wire12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_st_busy_wire130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_prot_true646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_wire23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range82w83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w661w806w807w817w818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode259w313w314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode259w260w261w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write86w87w442w443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_end_operation579w580w581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire446w447w448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy439w440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy431w432w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly600w601w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire476w477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire336w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode259w313w314w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode259w260w261w262w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w648w649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_rden_wire446w447w448w449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_not_busy431w432w433w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w263w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w316w317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w263w264w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w316w317w318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w263w264w265w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w316w317w318w319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w263w264w265w266w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w316w317w318w319w320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w263w264w265w266w267w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w316w317w318w319w320w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w263w264w265w266w267w268w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w269w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w322w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w269w270w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w322w323w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w269w270w271w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w322w323w324w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w269w270w271w272w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w322w323w324w325w326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w269w270w271w272w273w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w322w323w324w325w326w327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w269w270w271w272w273w274w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w275w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w328w329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w275w276w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w275w276w277w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w167w168w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w167w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w707w709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read335w462w463w464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read_sid163w164w165w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp3_wire670w671w672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read335w462w463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_sid163w164w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_stat342w343w344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_stat342w472w473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_erase663w664w665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write86w133w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_prot_wire_range683w701w703w705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp3_wire670w671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read335w475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read335w462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_rdid332w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_sid163w164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat346w347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat342w343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat342w472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase663w664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write86w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write86w87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly594w595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_prot_wire_range683w701w703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp3_wire670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data0out_wire479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_sid163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range720w748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range725w752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range730w756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range735w760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range739w764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range722w746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range727w750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range732w754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range737w758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range741w762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range612w615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range616w618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range619w621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range622w624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range625w627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range628w630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range631w633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range634w636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_prot_wire_range683w701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range699w715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range702w721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range704w726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range706w731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range708w736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range710w740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  add_rollover :	STD_LOGIC;
	 SIGNAL  addr_overdie :	STD_LOGIC;
	 SIGNAL  addr_overdie_pos :	STD_LOGIC;
	 SIGNAL  addr_reg_overdie :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  b4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  be_write_prot :	STD_LOGIC;
	 SIGNAL  berase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  bp0_wire :	STD_LOGIC;
	 SIGNAL  bp1_wire :	STD_LOGIC;
	 SIGNAL  bp2_wire :	STD_LOGIC;
	 SIGNAL  bp3_wire :	STD_LOGIC;
	 SIGNAL  buf_empty :	STD_LOGIC;
	 SIGNAL  busy_wire :	STD_LOGIC;
	 SIGNAL  clkin_wire :	STD_LOGIC;
	 SIGNAL  clr_addmsb_wire :	STD_LOGIC;
	 SIGNAL  clr_endrbyte_wire :	STD_LOGIC;
	 SIGNAL  clr_rdid_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire2 :	STD_LOGIC;
	 SIGNAL  clr_rstat_wire :	STD_LOGIC;
	 SIGNAL  clr_sid_wire :	STD_LOGIC;
	 SIGNAL  clr_write_wire :	STD_LOGIC;
	 SIGNAL  clr_write_wire2 :	STD_LOGIC;
	 SIGNAL  cnt_bfend_wire_in :	STD_LOGIC;
	 SIGNAL  data0out_wire :	STD_LOGIC;
	 SIGNAL  data_valid_wire :	STD_LOGIC;
	 SIGNAL  dataout_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  derase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  do_4baddr :	STD_LOGIC;
	 SIGNAL  do_bulk_erase :	STD_LOGIC;
	 SIGNAL  do_die_erase :	STD_LOGIC;
	 SIGNAL  do_ex4baddr :	STD_LOGIC;
	 SIGNAL  do_fast_read :	STD_LOGIC;
	 SIGNAL  do_fread_epcq :	STD_LOGIC;
	 SIGNAL  do_freadwrv_polling :	STD_LOGIC;
	 SIGNAL  do_memadd :	STD_LOGIC;
	 SIGNAL  do_polling :	STD_LOGIC;
	 SIGNAL  do_read :	STD_LOGIC;
	 SIGNAL  do_read_nonvolatile :	STD_LOGIC;
	 SIGNAL  do_read_rdid :	STD_LOGIC;
	 SIGNAL  do_read_sid :	STD_LOGIC;
	 SIGNAL  do_read_stat :	STD_LOGIC;
	 SIGNAL  do_read_volatile :	STD_LOGIC;
	 SIGNAL  do_sec_erase :	STD_LOGIC;
	 SIGNAL  do_sec_prot :	STD_LOGIC;
	 SIGNAL  do_secprot_wren :	STD_LOGIC;
	 SIGNAL  do_sprot_polling :	STD_LOGIC;
	 SIGNAL  do_sprot_rstat :	STD_LOGIC;
	 SIGNAL  do_wait_dummyclk :	STD_LOGIC;
	 SIGNAL  do_wren :	STD_LOGIC;
	 SIGNAL  do_write :	STD_LOGIC;
	 SIGNAL  do_write_polling :	STD_LOGIC;
	 SIGNAL  do_write_rstat :	STD_LOGIC;
	 SIGNAL  do_write_volatile :	STD_LOGIC;
	 SIGNAL  do_write_volatile_rstat :	STD_LOGIC;
	 SIGNAL  do_write_volatile_wren :	STD_LOGIC;
	 SIGNAL  do_write_wren :	STD_LOGIC;
	 SIGNAL  dummy_read_buf :	STD_LOGIC;
	 SIGNAL  end1_cyc_dlyncs_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_gen_cntr_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_normal_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_reg_in_wire :	STD_LOGIC;
	 SIGNAL  end_add_cycle :	STD_LOGIC;
	 SIGNAL  end_add_cycle_mux_datab_wire :	STD_LOGIC;
	 SIGNAL  end_fast_read :	STD_LOGIC;
	 SIGNAL  end_one_cyc_pos :	STD_LOGIC;
	 SIGNAL  end_one_cycle :	STD_LOGIC;
	 SIGNAL  end_op_wire :	STD_LOGIC;
	 SIGNAL  end_operation :	STD_LOGIC;
	 SIGNAL  end_ophdly :	STD_LOGIC;
	 SIGNAL  end_pgwr_data :	STD_LOGIC;
	 SIGNAL  end_read :	STD_LOGIC;
	 SIGNAL  end_read_byte :	STD_LOGIC;
	 SIGNAL  end_wrstage :	STD_LOGIC;
	 SIGNAL  exb4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fast_read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fast_read_wire :	STD_LOGIC;
	 SIGNAL  freadwrv_sdoin :	STD_LOGIC;
	 SIGNAL  ill_erase_wire :	STD_LOGIC;
	 SIGNAL  ill_write_wire :	STD_LOGIC;
	 SIGNAL  illegal_erase_b4out_wire :	STD_LOGIC;
	 SIGNAL  illegal_write_b4out_wire :	STD_LOGIC;
	 SIGNAL  in_operation :	STD_LOGIC;
	 SIGNAL  load_opcode :	STD_LOGIC;
	 SIGNAL  mask_prot :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mask_prot_add :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mask_prot_check :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mask_prot_comp_ntb :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mask_prot_comp_tb :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  memadd_sdoin :	STD_LOGIC;
	 SIGNAL  ncs_reg_ena_wire :	STD_LOGIC;
	 SIGNAL  not_busy :	STD_LOGIC;
	 SIGNAL  oe_wire :	STD_LOGIC;
	 SIGNAL  page_size_wire :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  pagewr_buf_not_empty :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  prot_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rden_wire :	STD_LOGIC;
	 SIGNAL  rdid_load :	STD_LOGIC;
	 SIGNAL  rdid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  reach_max_cnt :	STD_LOGIC;
	 SIGNAL  read_buf :	STD_LOGIC;
	 SIGNAL  read_bufdly :	STD_LOGIC;
	 SIGNAL  read_data_reg_in_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_rdid_wire :	STD_LOGIC;
	 SIGNAL  read_sid_wire :	STD_LOGIC;
	 SIGNAL  read_status_wire :	STD_LOGIC;
	 SIGNAL  read_wire :	STD_LOGIC;
	 SIGNAL  rflagstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rnvdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_sdoin :	STD_LOGIC;
	 SIGNAL  rstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  scein_wire :	STD_LOGIC;
	 SIGNAL  sdoin_wire :	STD_LOGIC;
	 SIGNAL  sec_erase_wire :	STD_LOGIC;
	 SIGNAL  sec_protect_wire :	STD_LOGIC;
	 SIGNAL  secprot_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  secprot_sdoin :	STD_LOGIC;
	 SIGNAL  serase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  shift_bytes_wire :	STD_LOGIC;
	 SIGNAL  shift_opcode :	STD_LOGIC;
	 SIGNAL  shift_opdata :	STD_LOGIC;
	 SIGNAL  shift_pgwr_data :	STD_LOGIC;
	 SIGNAL  st_busy_wire :	STD_LOGIC;
	 SIGNAL  stage2_wire :	STD_LOGIC;
	 SIGNAL  stage3_wire :	STD_LOGIC;
	 SIGNAL  stage4_wire :	STD_LOGIC;
	 SIGNAL  start_frpoll :	STD_LOGIC;
	 SIGNAL  start_poll :	STD_LOGIC;
	 SIGNAL  start_sppoll :	STD_LOGIC;
	 SIGNAL  start_wrpoll :	STD_LOGIC;
	 SIGNAL  to_sdoin_wire :	STD_LOGIC;
	 SIGNAL  wren_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wren_wire :	STD_LOGIC;
	 SIGNAL  write_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  write_prot_true :	STD_LOGIC;
	 SIGNAL  write_sdoin :	STD_LOGIC;
	 SIGNAL  write_wire :	STD_LOGIC;
	 SIGNAL  wrvolatile_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_addr_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_range430w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range426w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range191w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range199w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_dataout_wire_range478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range204w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_exb4addr_opcode_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exb4addr_opcode_range186w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range244w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range255w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range237w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range247w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range214w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range227w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range258w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range218w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range250w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range209w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range196w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range222w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range230w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 COMPONENT  a_graycounter
	 GENERIC 
	 (
		PVALUE	:	NATURAL := 0;
		WIDTH	:	NATURAL := 8;
		lpm_type	:	STRING := "a_graycounter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		q	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		qbin	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  scfifo
	 GENERIC 
	 (
		ADD_RAM_OUTPUT_REGISTER	:	STRING := "OFF";
		ALLOW_RWCYCLE_WHEN_FULL	:	STRING := "OFF";
		ALMOST_EMPTY_VALUE	:	NATURAL := 0;
		ALMOST_FULL_VALUE	:	NATURAL := 0;
		ENABLE_ECC	:	STRING := "FALSE";
		LPM_NUMWORDS	:	NATURAL;
		LPM_SHOWAHEAD	:	STRING := "OFF";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHU	:	NATURAL := 1;
		OVERFLOW_CHECKING	:	STRING := "ON";
		RAM_BLOCK_TYPE	:	STRING := "AUTO";
		UNDERFLOW_CHECKING	:	STRING := "ON";
		USE_EAB	:	STRING := "ON";
		lpm_type	:	STRING := "scfifo"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		almost_empty	:	OUT STD_LOGIC;
		almost_full	:	OUT STD_LOGIC;
		clock	:	IN STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		eccstatus	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		empty	:	OUT STD_LOGIC;
		full	:	OUT STD_LOGIC;
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		rdreq	:	IN STD_LOGIC;
		sclr	:	IN STD_LOGIC := '0';
		usedw	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHU-1 DOWNTO 0);
		wrreq	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_w568w569w570w571w(0) <= wire_w_lg_w_lg_w568w569w570w(0) AND wire_w_lg_do_ex4baddr557w(0);
	wire_w_lg_w_lg_w568w569w570w(0) <= wire_w_lg_w568w569w(0) AND wire_w_lg_do_4baddr558w(0);
	wire_w_lg_w_lg_w814w815w816w(0) <= wire_w_lg_w814w815w(0) AND end_operation;
	wire_w_lg_w568w569w(0) <= wire_w568w(0) AND wire_w_lg_do_sec_prot559w(0);
	wire_w_lg_w814w815w(0) <= wire_w814w(0) AND wire_w_lg_do_ex4baddr557w(0);
	wire_w568w(0) <= wire_w_lg_w_lg_w_lg_w_lg_end_ophdly564w565w566w567w(0) AND wire_w_lg_do_bulk_erase560w(0);
	wire_w303w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode239w240w241w242w(0) AND wire_w_rdummyclk_opcode_range302w(0);
	loop0 : FOR i IN 0 TO 6 GENERATE 
		wire_w243w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode239w240w241w242w(0) AND wire_w_rdummyclk_opcode_range237w(i);
	END GENERATE loop0;
	wire_w301w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode232w233w234w235w(0) AND wire_w_wrvolatile_opcode_range300w(0);
	loop1 : FOR i IN 0 TO 6 GENERATE 
		wire_w236w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode232w233w234w235w(0) AND wire_w_wrvolatile_opcode_range230w(i);
	END GENERATE loop1;
	wire_w814w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write563w811w812w813w(0) AND wire_w_lg_do_4baddr558w(0);
	wire_w510w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read335w507w508w509w(0) AND end_read_byte;
	wire_w_lg_w_lg_w_lg_w_lg_end_ophdly564w565w566w567w(0) <= wire_w_lg_w_lg_w_lg_end_ophdly564w565w566w(0) AND wire_w_lg_do_die_erase561w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode200w201w202w287w(0) <= wire_w_lg_w_lg_w_lg_load_opcode200w201w202w(0) AND wire_w_berase_opcode_range286w(0);
	loop2 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode200w201w202w203w(i) <= wire_w_lg_w_lg_w_lg_load_opcode200w201w202w(0) AND wire_w_berase_opcode_range199w(i);
	END GENERATE loop2;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w289w(0) <= wire_w_lg_w_lg_w_lg_load_opcode205w206w207w(0) AND wire_w_derase_opcode_range288w(0);
	loop3 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w(i) <= wire_w_lg_w_lg_w_lg_load_opcode205w206w207w(0) AND wire_w_derase_opcode_range204w(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode239w240w241w242w(0) <= wire_w_lg_w_lg_w_lg_load_opcode239w240w241w(0) AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode210w211w212w291w(0) <= wire_w_lg_w_lg_w_lg_load_opcode210w211w212w(0) AND wire_w_serase_opcode_range290w(0);
	loop4 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode210w211w212w213w(i) <= wire_w_lg_w_lg_w_lg_load_opcode210w211w212w(0) AND wire_w_serase_opcode_range209w(i);
	END GENERATE loop4;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode251w252w253w309w(0) <= wire_w_lg_w_lg_w_lg_load_opcode251w252w253w(0) AND wire_w_secprot_opcode_range308w(0);
	loop5 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode251w252w253w254w(i) <= wire_w_lg_w_lg_w_lg_load_opcode251w252w253w(0) AND wire_w_secprot_opcode_range250w(i);
	END GENERATE loop5;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode232w233w234w235w(0) <= wire_w_lg_w_lg_w_lg_load_opcode232w233w234w(0) AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_read394w395w396w397w(0) <= wire_w_lg_w_lg_w_lg_do_read394w395w396w(0) AND end_one_cycle;
	wire_w_lg_w_lg_w_lg_w_lg_do_write563w811w812w813w(0) <= wire_w_lg_w_lg_w_lg_do_write563w811w812w(0) AND wire_w_lg_do_die_erase561w(0);
	wire_w_lg_w_lg_w_lg_w661w806w807w817w(0) <= wire_w_lg_w_lg_w661w806w807w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_w_lg_do_read335w507w508w509w(0) <= wire_w_lg_w_lg_w_lg_do_read335w507w508w(0) AND end_one_cyc_pos;
	wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase68w450w451w452w(0) <= wire_w_lg_w_lg_w_lg_do_sec_erase68w450w451w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_end_ophdly564w565w566w(0) <= wire_w_lg_w_lg_end_ophdly564w565w(0) AND wire_w_lg_do_sec_erase562w(0);
	wire_w_lg_w_lg_w_lg_load_opcode200w201w202w(0) <= wire_w_lg_w_lg_load_opcode200w201w(0) AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_w_lg_w_lg_load_opcode205w206w207w(0) <= wire_w_lg_w_lg_load_opcode205w206w(0) AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_w_lg_w_lg_load_opcode215w220w295w(0) <= wire_w_lg_w_lg_load_opcode215w220w(0) AND wire_w_rstat_opcode_range294w(0);
	loop6 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode215w220w221w(i) <= wire_w_lg_w_lg_load_opcode215w220w(0) AND wire_w_rstat_opcode_range218w(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_w_lg_load_opcode215w216w293w(0) <= wire_w_lg_w_lg_load_opcode215w216w(0) AND wire_w_rflagstat_opcode_range292w(0);
	loop7 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode215w216w217w(i) <= wire_w_lg_w_lg_load_opcode215w216w(0) AND wire_w_rflagstat_opcode_range214w(i);
	END GENERATE loop7;
	wire_w_lg_w_lg_w_lg_load_opcode239w240w241w(0) <= wire_w_lg_w_lg_load_opcode239w240w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_w_lg_load_opcode210w211w212w(0) <= wire_w_lg_w_lg_load_opcode210w211w(0) AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_w_lg_w_lg_load_opcode251w252w253w(0) <= wire_w_lg_w_lg_load_opcode251w252w(0) AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_w_lg_w_lg_load_opcode232w233w234w(0) <= wire_w_lg_w_lg_load_opcode232w233w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_w_lg_bp2_wire677w678w679w(0) <= wire_w_lg_w_lg_bp2_wire677w678w(0) AND wire_w_lg_bp0_wire675w(0);
	wire_w_lg_w_lg_w_lg_bp2_wire677w678w682w(0) <= wire_w_lg_w_lg_bp2_wire677w678w(0) AND bp0_wire;
	wire_w_lg_w_lg_w_lg_bp2_wire677w684w685w(0) <= wire_w_lg_w_lg_bp2_wire677w684w(0) AND wire_w_lg_bp0_wire675w(0);
	wire_w_lg_w_lg_w_lg_bp2_wire677w684w687w(0) <= wire_w_lg_w_lg_bp2_wire677w684w(0) AND bp0_wire;
	wire_w_lg_w_lg_w_lg_do_read394w395w396w(0) <= wire_w_lg_w_lg_do_read394w395w(0) AND wire_w_lg_w_lg_do_write77w392w(0);
	wire_w_lg_w_lg_w_lg_do_read394w395w453w(0) <= wire_w_lg_w_lg_do_read394w395w(0) AND clr_write_wire2;
	wire_w_lg_w_lg_w_lg_do_write563w811w812w(0) <= wire_w_lg_w_lg_do_write563w811w(0) AND wire_w_lg_do_bulk_erase560w(0);
	wire_w_lg_w_lg_w661w806w807w(0) <= wire_w_lg_w661w806w(0) AND wire_wrstage_cntr_w_lg_w_q_range653w654w(0);
	wire_w_lg_w_lg_w_lg_do_read335w507w508w(0) <= wire_w_lg_w_lg_do_read335w507w(0) AND wire_stage_cntr_w_lg_w_q_range115w120w(0);
	wire_w_lg_w_lg_w_lg_do_sec_erase68w450w451w(0) <= wire_w_lg_w_lg_do_sec_erase68w450w(0) AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_w_lg_bp2_wire689w690w(0) <= wire_w_lg_bp2_wire689w(0) AND wire_w_lg_bp0_wire675w(0);
	wire_w_lg_w_lg_bp2_wire689w692w(0) <= wire_w_lg_bp2_wire689w(0) AND bp0_wire;
	wire_w_lg_w_lg_bp2_wire694w695w(0) <= wire_w_lg_bp2_wire694w(0) AND wire_w_lg_bp0_wire675w(0);
	wire_w_lg_w_lg_bp2_wire694w697w(0) <= wire_w_lg_bp2_wire694w(0) AND bp0_wire;
	wire_w_lg_w_lg_do_4baddr192w193w(0) <= wire_w_lg_do_4baddr192w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_do_ex4baddr187w188w(0) <= wire_w_lg_do_ex4baddr187w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_do_polling577w578w(0) <= wire_w_lg_do_polling577w(0) AND stage3_dly_reg;
	wire_w_lg_w_lg_do_write223w224w(0) <= wire_w_lg_do_write223w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_do_write77w373w(0) <= wire_w_lg_do_write77w(0) AND end_pgwr_data;
	wire_w_lg_w_lg_end_ophdly564w565w(0) <= wire_w_lg_end_ophdly564w(0) AND wire_w_lg_do_write563w(0);
	wire_w_lg_w_lg_end_read_byte514w526w(0) <= wire_w_lg_end_read_byte514w(0) AND wire_w_lg_end_operation525w(0);
	wire_w_lg_w_lg_load_opcode194w283w(0) <= wire_w_lg_load_opcode194w(0) AND wire_w_b4addr_opcode_range282w(0);
	loop8 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode194w195w(i) <= wire_w_lg_load_opcode194w(0) AND wire_w_b4addr_opcode_range191w(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_load_opcode189w281w(0) <= wire_w_lg_load_opcode189w(0) AND wire_w_exb4addr_opcode_range280w(0);
	loop9 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode189w190w(i) <= wire_w_lg_load_opcode189w(0) AND wire_w_exb4addr_opcode_range186w(i);
	END GENERATE loop9;
	wire_w_lg_w_lg_load_opcode225w297w(0) <= wire_w_lg_load_opcode225w(0) AND wire_w_write_opcode_range296w(0);
	loop10 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode225w226w(i) <= wire_w_lg_load_opcode225w(0) AND wire_w_write_opcode_range222w(i);
	END GENERATE loop10;
	wire_w_lg_w_lg_load_opcode200w201w(0) <= wire_w_lg_load_opcode200w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_load_opcode205w206w(0) <= wire_w_lg_load_opcode205w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_load_opcode245w305w(0) <= wire_w_lg_load_opcode245w(0) AND wire_w_fast_read_opcode_range304w(0);
	loop11 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode245w246w(i) <= wire_w_lg_load_opcode245w(0) AND wire_w_fast_read_opcode_range244w(i);
	END GENERATE loop11;
	wire_w_lg_w_lg_load_opcode248w307w(0) <= wire_w_lg_load_opcode248w(0) AND wire_w_read_opcode_range306w(0);
	loop12 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode248w249w(i) <= wire_w_lg_load_opcode248w(0) AND wire_w_read_opcode_range247w(i);
	END GENERATE loop12;
	wire_w_lg_w_lg_load_opcode228w299w(0) <= wire_w_lg_load_opcode228w(0) AND wire_w_rnvdummyclk_opcode_range298w(0);
	loop13 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode228w229w(i) <= wire_w_lg_load_opcode228w(0) AND wire_w_rnvdummyclk_opcode_range227w(i);
	END GENERATE loop13;
	wire_w_lg_w_lg_load_opcode256w311w(0) <= wire_w_lg_load_opcode256w(0) AND wire_w_rdid_opcode_range310w(0);
	loop14 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode256w257w(i) <= wire_w_lg_load_opcode256w(0) AND wire_w_rdid_opcode_range255w(i);
	END GENERATE loop14;
	wire_w_lg_w_lg_load_opcode259w313w(0) <= wire_w_lg_load_opcode259w(0) AND wire_w_rsid_opcode_range312w(0);
	loop15 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode259w260w(i) <= wire_w_lg_load_opcode259w(0) AND wire_w_rsid_opcode_range258w(i);
	END GENERATE loop15;
	wire_w_lg_w_lg_load_opcode215w220w(0) <= wire_w_lg_load_opcode215w(0) AND wire_w_lg_do_polling219w(0);
	wire_w_lg_w_lg_load_opcode215w216w(0) <= wire_w_lg_load_opcode215w(0) AND do_polling;
	wire_w_lg_w_lg_load_opcode239w240w(0) <= wire_w_lg_load_opcode239w(0) AND wire_w_lg_do_write_volatile238w(0);
	wire_w_lg_w_lg_load_opcode210w211w(0) <= wire_w_lg_load_opcode210w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_load_opcode251w252w(0) <= wire_w_lg_load_opcode251w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_load_opcode197w285w(0) <= wire_w_lg_load_opcode197w(0) AND wire_w_wren_opcode_range284w(0);
	loop16 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode197w198w(i) <= wire_w_lg_load_opcode197w(0) AND wire_w_wren_opcode_range196w(i);
	END GENERATE loop16;
	wire_w_lg_w_lg_load_opcode232w233w(0) <= wire_w_lg_load_opcode232w(0) AND wire_w_lg_do_read_volatile231w(0);
	wire_w_lg_w_lg_reach_max_cnt643w644w(0) <= wire_w_lg_reach_max_cnt643w(0) AND wren_wire;
	wire_w_lg_w_lg_stage3_wire59w60w(0) <= wire_w_lg_stage3_wire59w(0) AND do_wait_dummyclk;
	wire_w_lg_w_lg_start_poll380w381w(0) <= wire_w_lg_start_poll380w(0) AND do_polling;
	wire_w_lg_w_lg_bp2_wire677w678w(0) <= wire_w_lg_bp2_wire677w(0) AND wire_w_lg_bp1_wire676w(0);
	wire_w_lg_w_lg_bp2_wire677w684w(0) <= wire_w_lg_bp2_wire677w(0) AND bp1_wire;
	wire_w_lg_w_lg_do_read394w395w(0) <= wire_w_lg_do_read394w(0) AND wire_w_lg_do_fast_read393w(0);
	wire_w_lg_w_lg_do_write563w811w(0) <= wire_w_lg_do_write563w(0) AND wire_w_lg_do_sec_erase562w(0);
	loop17 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_read_bufdly597w598w(i) <= wire_w_lg_read_bufdly597w(0) AND wire_pgwrbuf_dataout_w_q_range596w(i);
	END GENERATE loop17;
	wire_w_lg_w_lg_w648w649w650w(0) <= wire_w_lg_w648w649w(0) AND end_wrstage;
	wire_w_lg_w661w806w(0) <= wire_w661w(0) AND wire_wrstage_cntr_w_q_range655w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w647w(0) <= wire_w_lg_w_lg_w_lg_do_write86w133w134w(0) AND wire_w_lg_write_prot_true646w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w135w(0) <= wire_w_lg_w_lg_w_lg_do_write86w133w134w(0) AND write_prot_true;
	wire_w_lg_w_lg_w_lg_do_write86w87w442w(0) <= wire_w_lg_w_lg_do_write86w87w(0) AND do_memadd;
	wire_w_lg_w_lg_do_read335w507w(0) <= wire_w_lg_do_read335w(0) AND wire_stage_cntr_w_q_range116w(0);
	wire_w_lg_w_lg_do_sec_erase68w450w(0) <= wire_w_lg_do_sec_erase68w(0) AND wire_w_lg_do_wren67w(0);
	wire_w_lg_w_lg_end_operation579w580w(0) <= wire_w_lg_end_operation579w(0) AND do_read_stat;
	wire_w_lg_w_lg_rden_wire446w447w(0) <= wire_w_lg_rden_wire446w(0) AND not_busy;
	wire_w_lg_addr_overdie437w(0) <= addr_overdie AND wire_w_addr_reg_overdie_range436w(0);
	loop18 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_addr_overdie427w(i) <= addr_overdie AND wire_w_addr_reg_overdie_range426w(i);
	END GENERATE loop18;
	wire_w_lg_bp2_wire689w(0) <= bp2_wire AND wire_w_lg_bp1_wire676w(0);
	wire_w_lg_bp2_wire694w(0) <= bp2_wire AND bp1_wire;
	wire_w_lg_do_4baddr192w(0) <= do_4baddr AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_do_bulk_erase374w(0) <= do_bulk_erase AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_do_ex4baddr187w(0) <= do_ex4baddr AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_do_polling577w(0) <= do_polling AND end_one_cyc_pos;
	wire_w_lg_do_read_nonvolatile360w(0) <= do_read_nonvolatile AND wire_addbyte_cntr_w_q_range174w(0);
	wire_w_lg_do_write223w(0) <= do_write AND wire_w_lg_do_read_stat66w(0);
	wire_w_lg_do_write84w(0) <= do_write AND wire_w_lg_w_pagewr_buf_not_empty_range82w83w(0);
	wire_w_lg_do_write77w(0) <= do_write AND shift_pgwr_data;
	wire_w_lg_end_operation545w(0) <= end_operation AND wire_w_lg_do_read335w(0);
	wire_w_lg_end_ophdly564w(0) <= end_ophdly AND do_read_stat;
	wire_w_lg_end_read_byte514w(0) <= end_read_byte AND end_one_cyc_pos;
	wire_w_lg_in_operation52w(0) <= in_operation AND wire_w_lg_end_ophdly51w(0);
	wire_w_lg_load_opcode194w(0) <= load_opcode AND wire_w_lg_w_lg_do_4baddr192w193w(0);
	wire_w_lg_load_opcode189w(0) <= load_opcode AND wire_w_lg_w_lg_do_ex4baddr187w188w(0);
	wire_w_lg_load_opcode225w(0) <= load_opcode AND wire_w_lg_w_lg_do_write223w224w(0);
	wire_w_lg_load_opcode200w(0) <= load_opcode AND do_bulk_erase;
	wire_w_lg_load_opcode205w(0) <= load_opcode AND do_die_erase;
	wire_w_lg_load_opcode245w(0) <= load_opcode AND do_fast_read;
	wire_w_lg_load_opcode248w(0) <= load_opcode AND do_read;
	wire_w_lg_load_opcode228w(0) <= load_opcode AND do_read_nonvolatile;
	wire_w_lg_load_opcode256w(0) <= load_opcode AND do_read_rdid;
	wire_w_lg_load_opcode259w(0) <= load_opcode AND do_read_sid;
	wire_w_lg_load_opcode215w(0) <= load_opcode AND do_read_stat;
	wire_w_lg_load_opcode239w(0) <= load_opcode AND do_read_volatile;
	wire_w_lg_load_opcode210w(0) <= load_opcode AND do_sec_erase;
	wire_w_lg_load_opcode251w(0) <= load_opcode AND do_sec_prot;
	wire_w_lg_load_opcode197w(0) <= load_opcode AND do_wren;
	wire_w_lg_load_opcode232w(0) <= load_opcode AND do_write_volatile;
	wire_w_lg_not_busy439w(0) <= not_busy AND wire_w_addr_range438w(0);
	loop19 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_not_busy431w(i) <= not_busy AND wire_w_addr_range430w(i);
	END GENERATE loop19;
	wire_w_lg_reach_max_cnt643w(0) <= reach_max_cnt AND shift_bytes_wire;
	wire_w_lg_read_bufdly605w(0) <= read_bufdly AND wire_scfifo3_w_q_range604w(0);
	loop20 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_read_bufdly600w(i) <= read_bufdly AND wire_scfifo3_w_q_range599w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_shift_opcode185w(i) <= shift_opcode AND wire_asmi_opcode_reg_w_q_range184w(i);
	END GENERATE loop21;
	wire_w_lg_stage3_wire444w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_w_lg_do_write86w87w442w443w(0);
	wire_w_lg_stage3_wire345w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_do_read_stat342w343w344w(0);
	wire_w_lg_stage3_wire474w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_do_read_stat342w472w473w(0);
	wire_w_lg_stage3_wire334w(0) <= stage3_wire AND wire_w_lg_w_lg_do_read_rdid332w333w(0);
	wire_w_lg_stage3_wire69w(0) <= stage3_wire AND wire_w_lg_do_sec_erase68w(0);
	wire_w_lg_stage3_wire59w(0) <= stage3_wire AND do_fast_read;
	loop22 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_stage3_wire429w(i) <= stage3_wire AND wire_addr_reg_w_q_range428w(i);
	END GENERATE loop22;
	wire_w_lg_stage4_wire476w(0) <= stage4_wire AND wire_w_lg_w_lg_do_read335w475w(0);
	wire_w_lg_stage4_wire336w(0) <= stage4_wire AND wire_w_lg_do_read335w(0);
	wire_w_lg_stage4_wire445w(0) <= stage4_wire AND addr_overdie;
	wire_w_lg_stage4_wire350w(0) <= stage4_wire AND do_fast_read;
	wire_w_lg_start_poll380w(0) <= start_poll AND do_read_stat;
	wire_w_lg_w_mask_prot_range699w712w(0) <= wire_w_mask_prot_range699w(0) AND wire_addr_reg_w_q_range711w(0);
	wire_w_lg_w_mask_prot_range702w719w(0) <= wire_w_mask_prot_range702w(0) AND wire_addr_reg_w_q_range718w(0);
	wire_w_lg_w_mask_prot_range704w724w(0) <= wire_w_mask_prot_range704w(0) AND wire_addr_reg_w_q_range723w(0);
	wire_w_lg_w_mask_prot_range706w729w(0) <= wire_w_mask_prot_range706w(0) AND wire_addr_reg_w_q_range728w(0);
	wire_w_lg_w_mask_prot_range708w734w(0) <= wire_w_mask_prot_range708w(0) AND wire_addr_reg_w_q_range733w(0);
	wire_w_lg_w_mask_prot_range710w738w(0) <= wire_w_mask_prot_range710w(0) AND wire_addr_reg_w_q_range458w(0);
	wire_w_lg_w_lg_do_write77w392w(0) <= NOT wire_w_lg_do_write77w(0);
	wire_w_lg_w_lg_stage4_wire350w351w(0) <= NOT wire_w_lg_stage4_wire350w(0);
	wire_w_lg_w_lg_w_lg_stage4_wire336w337w338w(0) <= NOT wire_w_lg_w_lg_stage4_wire336w337w(0);
	wire_w_lg_w_lg_w_lg_do_read_stat346w347w348w(0) <= NOT wire_w_lg_w_lg_do_read_stat346w347w(0);
	wire_w_lg_addr_overdie539w(0) <= NOT addr_overdie;
	wire_w_lg_bp0_wire675w(0) <= NOT bp0_wire;
	wire_w_lg_bp1_wire676w(0) <= NOT bp1_wire;
	wire_w_lg_bp2_wire677w(0) <= NOT bp2_wire;
	wire_w_lg_buf_empty780w(0) <= NOT buf_empty;
	wire_w_lg_busy_wire3w(0) <= NOT busy_wire;
	wire_w_lg_clkin_wire48w(0) <= NOT clkin_wire;
	wire_w_lg_clr_rstat_wire50w(0) <= NOT clr_rstat_wire;
	wire_w_lg_clr_sid_wire49w(0) <= NOT clr_sid_wire;
	wire_w_lg_do_4baddr558w(0) <= NOT do_4baddr;
	wire_w_lg_do_bulk_erase560w(0) <= NOT do_bulk_erase;
	wire_w_lg_do_die_erase561w(0) <= NOT do_die_erase;
	wire_w_lg_do_ex4baddr557w(0) <= NOT do_ex4baddr;
	wire_w_lg_do_fast_read393w(0) <= NOT do_fast_read;
	wire_w_lg_do_memadd459w(0) <= NOT do_memadd;
	wire_w_lg_do_polling219w(0) <= NOT do_polling;
	wire_w_lg_do_read394w(0) <= NOT do_read;
	wire_w_lg_do_read_nonvolatile10w(0) <= NOT do_read_nonvolatile;
	wire_w_lg_do_read_rdid65w(0) <= NOT do_read_rdid;
	wire_w_lg_do_read_stat66w(0) <= NOT do_read_stat;
	wire_w_lg_do_read_volatile231w(0) <= NOT do_read_volatile;
	wire_w_lg_do_sec_erase562w(0) <= NOT do_sec_erase;
	wire_w_lg_do_sec_prot559w(0) <= NOT do_sec_prot;
	wire_w_lg_do_wren67w(0) <= NOT do_wren;
	wire_w_lg_do_write563w(0) <= NOT do_write;
	wire_w_lg_do_write_volatile238w(0) <= NOT do_write_volatile;
	wire_w_lg_end_add_cycle97w(0) <= NOT end_add_cycle;
	wire_w_lg_end_fast_read91w(0) <= NOT end_fast_read;
	wire_w_lg_end_operation525w(0) <= NOT end_operation;
	wire_w_lg_end_ophdly51w(0) <= NOT end_ophdly;
	wire_w_lg_end_pgwr_data76w(0) <= NOT end_pgwr_data;
	wire_w_lg_end_read94w(0) <= NOT end_read;
	wire_w_lg_rden_wire541w(0) <= NOT rden_wire;
	wire_w_lg_reach_max_cnt607w(0) <= NOT reach_max_cnt;
	wire_w_lg_read_bufdly597w(0) <= NOT read_bufdly;
	wire_w_lg_read_rdid_wire14w(0) <= NOT read_rdid_wire;
	wire_w_lg_read_sid_wire13w(0) <= NOT read_sid_wire;
	wire_w_lg_read_status_wire29w(0) <= NOT read_status_wire;
	wire_w_lg_sec_protect_wire12w(0) <= NOT sec_protect_wire;
	wire_w_lg_st_busy_wire130w(0) <= NOT st_busy_wire;
	wire_w_lg_write_prot_true646w(0) <= NOT write_prot_true;
	wire_w_lg_write_wire23w(0) <= NOT write_wire;
	wire_w_lg_w_pagewr_buf_not_empty_range82w83w(0) <= NOT wire_w_pagewr_buf_not_empty_range82w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w661w806w807w817w818w(0) <= wire_w_lg_w_lg_w_lg_w661w806w807w817w(0) OR write_prot_true;
	wire_w_lg_w_lg_w_lg_load_opcode259w313w314w(0) <= wire_w_lg_w_lg_load_opcode259w313w(0) OR wire_w_lg_w_lg_load_opcode256w311w(0);
	loop23 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode259w260w261w(i) <= wire_w_lg_w_lg_load_opcode259w260w(i) OR wire_w_lg_w_lg_load_opcode256w257w(i);
	END GENERATE loop23;
	wire_w648w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w647w(0) OR do_4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_do_write86w87w442w443w(0) <= wire_w_lg_w_lg_w_lg_do_write86w87w442w(0) OR wire_w_lg_do_read335w(0);
	wire_w_lg_w_lg_w_lg_end_operation579w580w581w(0) <= wire_w_lg_w_lg_end_operation579w580w(0) OR clr_rstat_wire;
	wire_w_lg_w_lg_w_lg_rden_wire446w447w448w(0) <= wire_w_lg_w_lg_rden_wire446w447w(0) OR wire_w_lg_stage4_wire445w(0);
	wire_w_lg_w_lg_not_busy439w440w(0) <= wire_w_lg_not_busy439w(0) OR wire_w_lg_addr_overdie437w(0);
	loop24 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_not_busy431w432w(i) <= wire_w_lg_not_busy431w(i) OR wire_w_lg_stage3_wire429w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_read_bufdly600w601w(i) <= wire_w_lg_read_bufdly600w(i) OR wire_w_lg_w_lg_read_bufdly597w598w(i);
	END GENERATE loop25;
	wire_w_lg_w_lg_stage4_wire476w477w(0) <= wire_w_lg_stage4_wire476w(0) OR wire_w_lg_stage3_wire474w(0);
	wire_w_lg_w_lg_stage4_wire336w337w(0) <= wire_w_lg_stage4_wire336w(0) OR wire_w_lg_stage3_wire334w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode259w313w314w315w(0) <= wire_w_lg_w_lg_w_lg_load_opcode259w313w314w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode251w252w253w309w(0);
	loop26 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode259w260w261w262w(i) <= wire_w_lg_w_lg_w_lg_load_opcode259w260w261w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode251w252w253w254w(i);
	END GENERATE loop26;
	wire_w_lg_w648w649w(0) <= wire_w648w(0) OR do_ex4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_rden_wire446w447w448w449w(0) <= wire_w_lg_w_lg_w_lg_rden_wire446w447w448w(0) OR wire_w_lg_stage3_wire444w(0);
	loop27 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_w_lg_not_busy431w432w433w(i) <= wire_w_lg_w_lg_not_busy431w432w(i) OR wire_w_lg_addr_overdie427w(i);
	END GENERATE loop27;
	wire_w316w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode259w313w314w315w(0) OR wire_w_lg_w_lg_load_opcode248w307w(0);
	loop28 : FOR i IN 0 TO 6 GENERATE 
		wire_w263w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode259w260w261w262w(i) OR wire_w_lg_w_lg_load_opcode248w249w(i);
	END GENERATE loop28;
	wire_w_lg_w316w317w(0) <= wire_w316w(0) OR wire_w_lg_w_lg_load_opcode245w305w(0);
	loop29 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w263w264w(i) <= wire_w263w(i) OR wire_w_lg_w_lg_load_opcode245w246w(i);
	END GENERATE loop29;
	wire_w_lg_w_lg_w316w317w318w(0) <= wire_w_lg_w316w317w(0) OR wire_w303w(0);
	loop30 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w263w264w265w(i) <= wire_w_lg_w263w264w(i) OR wire_w243w(i);
	END GENERATE loop30;
	wire_w_lg_w_lg_w_lg_w316w317w318w319w(0) <= wire_w_lg_w_lg_w316w317w318w(0) OR wire_w301w(0);
	loop31 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w263w264w265w266w(i) <= wire_w_lg_w_lg_w263w264w265w(i) OR wire_w236w(i);
	END GENERATE loop31;
	wire_w_lg_w_lg_w_lg_w_lg_w316w317w318w319w320w(0) <= wire_w_lg_w_lg_w_lg_w316w317w318w319w(0) OR wire_w_lg_w_lg_load_opcode228w299w(0);
	loop32 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w263w264w265w266w267w(i) <= wire_w_lg_w_lg_w_lg_w263w264w265w266w(i) OR wire_w_lg_w_lg_load_opcode228w229w(i);
	END GENERATE loop32;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w316w317w318w319w320w321w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w316w317w318w319w320w(0) OR wire_w_lg_w_lg_load_opcode225w297w(0);
	loop33 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w263w264w265w266w267w268w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w263w264w265w266w267w(i) OR wire_w_lg_w_lg_load_opcode225w226w(i);
	END GENERATE loop33;
	wire_w322w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w316w317w318w319w320w321w(0) OR wire_w_lg_w_lg_w_lg_load_opcode215w220w295w(0);
	loop34 : FOR i IN 0 TO 6 GENERATE 
		wire_w269w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w263w264w265w266w267w268w(i) OR wire_w_lg_w_lg_w_lg_load_opcode215w220w221w(i);
	END GENERATE loop34;
	wire_w_lg_w322w323w(0) <= wire_w322w(0) OR wire_w_lg_w_lg_w_lg_load_opcode215w216w293w(0);
	loop35 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w269w270w(i) <= wire_w269w(i) OR wire_w_lg_w_lg_w_lg_load_opcode215w216w217w(i);
	END GENERATE loop35;
	wire_w_lg_w_lg_w322w323w324w(0) <= wire_w_lg_w322w323w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode210w211w212w291w(0);
	loop36 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w269w270w271w(i) <= wire_w_lg_w269w270w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode210w211w212w213w(i);
	END GENERATE loop36;
	wire_w_lg_w_lg_w_lg_w322w323w324w325w(0) <= wire_w_lg_w_lg_w322w323w324w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w289w(0);
	loop37 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w269w270w271w272w(i) <= wire_w_lg_w_lg_w269w270w271w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w(i);
	END GENERATE loop37;
	wire_w_lg_w_lg_w_lg_w_lg_w322w323w324w325w326w(0) <= wire_w_lg_w_lg_w_lg_w322w323w324w325w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode200w201w202w287w(0);
	loop38 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w269w270w271w272w273w(i) <= wire_w_lg_w_lg_w_lg_w269w270w271w272w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode200w201w202w203w(i);
	END GENERATE loop38;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w322w323w324w325w326w327w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w322w323w324w325w326w(0) OR wire_w_lg_w_lg_load_opcode197w285w(0);
	loop39 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w269w270w271w272w273w274w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w269w270w271w272w273w(i) OR wire_w_lg_w_lg_load_opcode197w198w(i);
	END GENERATE loop39;
	wire_w328w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w322w323w324w325w326w327w(0) OR wire_w_lg_w_lg_load_opcode194w283w(0);
	loop40 : FOR i IN 0 TO 6 GENERATE 
		wire_w275w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w269w270w271w272w273w274w(i) OR wire_w_lg_w_lg_load_opcode194w195w(i);
	END GENERATE loop40;
	wire_w_lg_w328w329w(0) <= wire_w328w(0) OR wire_w_lg_w_lg_load_opcode189w281w(0);
	loop41 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w275w276w(i) <= wire_w275w(i) OR wire_w_lg_w_lg_load_opcode189w190w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w275w276w277w(i) <= wire_w_lg_w275w276w(i) OR wire_w_lg_shift_opcode185w(i);
	END GENERATE loop42;
	wire_w_lg_w_lg_w167w168w169w(0) <= wire_w_lg_w167w168w(0) OR do_read_nonvolatile;
	wire_w_lg_w167w168w(0) <= wire_w167w(0) OR do_fast_read;
	wire_w167w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read_sid163w164w165w166w(0) OR do_read;
	wire_w661w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w660w(0) OR do_ex4baddr;
	wire_w_lg_w707w709w(0) <= wire_w707w(0) OR wire_w_prot_wire_range696w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_read335w462w463w464w(0) <= wire_w_lg_w_lg_w_lg_do_read335w462w463w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_w_lg_do_read_sid163w164w165w166w(0) <= wire_w_lg_w_lg_w_lg_do_read_sid163w164w165w(0) OR do_read_rdid;
	wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w660w(0) <= wire_w_lg_w_lg_w_lg_do_write86w133w134w(0) OR do_4baddr;
	wire_w707w(0) <= wire_w_lg_w_lg_w_lg_w_prot_wire_range683w701w703w705w(0) OR wire_w_prot_wire_range693w(0);
	wire_w_lg_w_lg_w_lg_bp3_wire670w671w672w(0) <= wire_w_lg_w_lg_bp3_wire670w671w(0) OR bp0_wire;
	wire_w_lg_w_lg_w_lg_do_read335w462w463w(0) <= wire_w_lg_w_lg_do_read335w462w(0) OR do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read_sid163w164w165w(0) <= wire_w_lg_w_lg_do_read_sid163w164w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_do_read_stat342w343w344w(0) <= wire_w_lg_w_lg_do_read_stat342w343w(0) OR do_read_volatile;
	wire_w_lg_w_lg_w_lg_do_read_stat342w472w473w(0) <= wire_w_lg_w_lg_do_read_stat342w472w(0) OR do_read_nonvolatile;
	wire_w_lg_w_lg_w_lg_do_sec_erase663w664w665w(0) <= wire_w_lg_w_lg_do_sec_erase663w664w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_do_write86w133w134w(0) <= wire_w_lg_w_lg_do_write86w133w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_w_prot_wire_range683w701w703w705w(0) <= wire_w_lg_w_lg_w_prot_wire_range683w701w703w(0) OR wire_w_prot_wire_range691w(0);
	wire_w_lg_w_lg_bp3_wire670w671w(0) <= wire_w_lg_bp3_wire670w(0) OR bp1_wire;
	wire_w_lg_w_lg_do_read335w475w(0) <= wire_w_lg_do_read335w(0) OR do_read_sid;
	wire_w_lg_w_lg_do_read335w462w(0) <= wire_w_lg_do_read335w(0) OR do_write;
	wire_w_lg_w_lg_do_read_rdid332w333w(0) <= wire_w_lg_do_read_rdid332w(0) OR do_read_volatile;
	wire_w_lg_w_lg_do_read_sid163w164w(0) <= wire_w_lg_do_read_sid163w(0) OR do_sec_erase;
	wire_w_lg_w_lg_do_read_stat346w347w(0) <= wire_w_lg_do_read_stat346w(0) OR wire_w_lg_stage3_wire345w(0);
	wire_w_lg_w_lg_do_read_stat342w343w(0) <= wire_w_lg_do_read_stat342w(0) OR do_read_nonvolatile;
	wire_w_lg_w_lg_do_read_stat342w472w(0) <= wire_w_lg_do_read_stat342w(0) OR do_read_volatile;
	wire_w_lg_w_lg_do_sec_erase663w664w(0) <= wire_w_lg_do_sec_erase663w(0) OR do_bulk_erase;
	wire_w_lg_w_lg_do_write86w133w(0) <= wire_w_lg_do_write86w(0) OR do_bulk_erase;
	wire_w_lg_w_lg_do_write86w87w(0) <= wire_w_lg_do_write86w(0) OR do_die_erase;
	wire_w_lg_w_lg_read_bufdly594w595w(0) <= wire_w_lg_read_bufdly594w(0) OR clr_write_wire;
	wire_w_lg_w_lg_w_prot_wire_range683w701w703w(0) <= wire_w_lg_w_prot_wire_range683w701w(0) OR wire_w_prot_wire_range688w(0);
	wire_w_lg_bp3_wire670w(0) <= bp3_wire OR bp2_wire;
	wire_w_lg_data0out_wire479w(0) <= data0out_wire OR wire_w_dataout_wire_range478w(0);
	wire_w_lg_do_4baddr376w(0) <= do_4baddr OR wire_w_lg_do_ex4baddr375w(0);
	wire_w_lg_do_ex4baddr375w(0) <= do_ex4baddr OR wire_w_lg_do_bulk_erase374w(0);
	wire_w_lg_do_read335w(0) <= do_read OR do_fast_read;
	wire_w_lg_do_read_rdid332w(0) <= do_read_rdid OR do_read_nonvolatile;
	wire_w_lg_do_read_sid163w(0) <= do_read_sid OR do_write;
	wire_w_lg_do_read_stat346w(0) <= do_read_stat OR wire_w_lg_stage4_wire336w(0);
	wire_w_lg_do_read_stat339w(0) <= do_read_stat OR wire_w_lg_w_lg_w_lg_stage4_wire336w337w338w(0);
	wire_w_lg_do_read_stat342w(0) <= do_read_stat OR do_read_rdid;
	wire_w_lg_do_sec_erase68w(0) <= do_sec_erase OR do_die_erase;
	wire_w_lg_do_sec_erase663w(0) <= do_sec_erase OR do_write;
	wire_w_lg_do_wren377w(0) <= do_wren OR wire_w_lg_do_4baddr376w(0);
	wire_w_lg_do_write86w(0) <= do_write OR do_sec_erase;
	wire_w_lg_end_operation579w(0) <= end_operation OR wire_w_lg_w_lg_do_polling577w578w(0);
	wire_w_lg_load_opcode331w(0) <= load_opcode OR shift_opcode;
	wire_w_lg_rden_wire446w(0) <= rden_wire OR wren_wire;
	wire_w_lg_read_bufdly594w(0) <= read_bufdly OR shift_pgwr_data;
	wire_w_lg_w_mask_prot_add_range720w748w(0) <= wire_w_mask_prot_add_range720w(0) OR wire_w_mask_prot_comp_tb_range744w(0);
	wire_w_lg_w_mask_prot_add_range725w752w(0) <= wire_w_mask_prot_add_range725w(0) OR wire_w_mask_prot_comp_tb_range749w(0);
	wire_w_lg_w_mask_prot_add_range730w756w(0) <= wire_w_mask_prot_add_range730w(0) OR wire_w_mask_prot_comp_tb_range753w(0);
	wire_w_lg_w_mask_prot_add_range735w760w(0) <= wire_w_mask_prot_add_range735w(0) OR wire_w_mask_prot_comp_tb_range757w(0);
	wire_w_lg_w_mask_prot_add_range739w764w(0) <= wire_w_mask_prot_add_range739w(0) OR wire_w_mask_prot_comp_tb_range761w(0);
	wire_w_lg_w_mask_prot_check_range722w746w(0) <= wire_w_mask_prot_check_range722w(0) OR wire_w_mask_prot_comp_ntb_range742w(0);
	wire_w_lg_w_mask_prot_check_range727w750w(0) <= wire_w_mask_prot_check_range727w(0) OR wire_w_mask_prot_comp_ntb_range747w(0);
	wire_w_lg_w_mask_prot_check_range732w754w(0) <= wire_w_mask_prot_check_range732w(0) OR wire_w_mask_prot_comp_ntb_range751w(0);
	wire_w_lg_w_mask_prot_check_range737w758w(0) <= wire_w_mask_prot_check_range737w(0) OR wire_w_mask_prot_comp_ntb_range755w(0);
	wire_w_lg_w_mask_prot_check_range741w762w(0) <= wire_w_mask_prot_check_range741w(0) OR wire_w_mask_prot_comp_ntb_range759w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range612w615w(0) <= wire_w_pagewr_buf_not_empty_range612w(0) OR wire_pgwr_data_cntr_w_q_range614w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range616w618w(0) <= wire_w_pagewr_buf_not_empty_range616w(0) OR wire_pgwr_data_cntr_w_q_range617w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range619w621w(0) <= wire_w_pagewr_buf_not_empty_range619w(0) OR wire_pgwr_data_cntr_w_q_range620w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range622w624w(0) <= wire_w_pagewr_buf_not_empty_range622w(0) OR wire_pgwr_data_cntr_w_q_range623w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range625w627w(0) <= wire_w_pagewr_buf_not_empty_range625w(0) OR wire_pgwr_data_cntr_w_q_range626w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range628w630w(0) <= wire_w_pagewr_buf_not_empty_range628w(0) OR wire_pgwr_data_cntr_w_q_range629w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range631w633w(0) <= wire_w_pagewr_buf_not_empty_range631w(0) OR wire_pgwr_data_cntr_w_q_range632w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range634w636w(0) <= wire_w_pagewr_buf_not_empty_range634w(0) OR wire_pgwr_data_cntr_w_q_range635w(0);
	wire_w_lg_w_prot_wire_range683w701w(0) <= wire_w_prot_wire_range683w(0) OR wire_w_prot_wire_range686w(0);
	wire_w_lg_w_mask_prot_range699w715w(0) <= wire_w_mask_prot_range699w(0) XOR wire_w_mask_prot_add_range713w(0);
	wire_w_lg_w_mask_prot_range702w721w(0) <= wire_w_mask_prot_range702w(0) XOR wire_w_mask_prot_add_range720w(0);
	wire_w_lg_w_mask_prot_range704w726w(0) <= wire_w_mask_prot_range704w(0) XOR wire_w_mask_prot_add_range725w(0);
	wire_w_lg_w_mask_prot_range706w731w(0) <= wire_w_mask_prot_range706w(0) XOR wire_w_mask_prot_add_range730w(0);
	wire_w_lg_w_mask_prot_range708w736w(0) <= wire_w_mask_prot_range708w(0) XOR wire_w_mask_prot_add_range735w(0);
	wire_w_lg_w_mask_prot_range710w740w(0) <= wire_w_mask_prot_range710w(0) XOR wire_w_mask_prot_add_range739w(0);
	add_rollover <= add_rollover_reg;
	addr_overdie <= '0';
	addr_overdie_pos <= '0';
	addr_reg_overdie <= (OTHERS => '0');
	asmi_dataoe <= oe_wire;
	asmi_dclk <= clkin_wire;
	asmi_scein <= scein_wire;
	asmi_sdoin <= sdoin_wire;
	b4addr_opcode <= (OTHERS => '0');
	be_write_prot <= ((do_bulk_erase OR do_die_erase) AND wire_w_lg_w_lg_w_lg_bp3_wire670w671w672w(0));
	berase_opcode <= (OTHERS => '0');
	bp0_wire <= statreg_int(2);
	bp1_wire <= statreg_int(3);
	bp2_wire <= statreg_int(4);
	bp3_wire <= statreg_int(6);
	buf_empty <= buf_empty_reg;
	busy <= (busy_wire OR busy_delay_reg);
	busy_wire <= ((((((((((((((do_read_rdid OR do_read_sid) OR do_read) OR do_fast_read) OR do_write) OR do_sec_prot) OR do_read_stat) OR do_sec_erase) OR do_bulk_erase) OR do_die_erase) OR do_4baddr) OR do_read_volatile) OR do_fread_epcq) OR do_read_nonvolatile) OR do_ex4baddr);
	clkin_wire <= clkin;
	clr_addmsb_wire <= ((wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w121w454w455w(0) OR wire_w_lg_w_lg_w_lg_do_read394w395w453w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase68w450w451w452w(0));
	clr_endrbyte_wire <= ((((wire_w_lg_do_read335w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR clr_read_wire2);
	clr_rdid_wire <= clr_rdid_reg;
	clr_read_wire <= clr_read_reg;
	clr_read_wire2 <= clr_read_reg2;
	clr_rstat_wire <= clr_rstat_reg;
	clr_sid_wire <= '0';
	clr_write_wire <= clr_write_reg;
	clr_write_wire2 <= clr_write_reg2;
	cnt_bfend_wire_in <= (wire_gen_cntr_w_lg_w_q_range126w127w(0) AND wire_gen_cntr_q(0));
	data0out_wire <= asmi_dataout;
	data_valid <= data_valid_wire;
	data_valid_wire <= dvalid_reg2;
	dataout <= ( read_data_reg(7 DOWNTO 0));
	dataout_wire <= ( "0000");
	derase_opcode <= (OTHERS => '0');
	do_4baddr <= '0';
	do_bulk_erase <= '0';
	do_die_erase <= '0';
	do_ex4baddr <= '0';
	do_fast_read <= ((((wire_w_lg_do_read_nonvolatile10w(0) AND wire_w_lg_read_rdid_wire14w(0)) AND wire_w_lg_read_sid_wire13w(0)) AND wire_w_lg_sec_protect_wire12w(0)) AND fast_read_wire);
	do_fread_epcq <= '0';
	do_freadwrv_polling <= '0';
	do_memadd <= do_wrmemadd_reg;
	do_polling <= ((do_write_polling OR do_sprot_polling) OR do_freadwrv_polling);
	do_read <= '0';
	do_read_nonvolatile <= '0';
	do_read_rdid <= (wire_w_lg_do_read_nonvolatile10w(0) AND read_rdid_wire);
	do_read_sid <= '0';
	do_read_stat <= (((((((((wire_w_lg_do_read_nonvolatile10w(0) AND wire_w_lg_read_rdid_wire14w(0)) AND wire_w_lg_read_sid_wire13w(0)) AND wire_w_lg_sec_protect_wire12w(0)) AND (NOT (read_wire OR fast_read_wire))) AND wire_w_lg_write_wire23w(0)) AND read_status_wire) OR do_write_rstat) OR do_sprot_rstat) OR do_write_volatile_rstat);
	do_read_volatile <= '0';
	do_sec_erase <= (((((((wire_w_lg_do_read_nonvolatile10w(0) AND wire_w_lg_read_rdid_wire14w(0)) AND wire_w_lg_read_sid_wire13w(0)) AND wire_w_lg_sec_protect_wire12w(0)) AND (NOT (read_wire OR fast_read_wire))) AND wire_w_lg_write_wire23w(0)) AND wire_w_lg_read_status_wire29w(0)) AND sec_erase_wire);
	do_sec_prot <= '0';
	do_secprot_wren <= '0';
	do_sprot_polling <= '0';
	do_sprot_rstat <= '0';
	do_wait_dummyclk <= '0';
	do_wren <= ((do_write_wren OR do_secprot_wren) OR do_write_volatile_wren);
	do_write <= (((((wire_w_lg_do_read_nonvolatile10w(0) AND wire_w_lg_read_rdid_wire14w(0)) AND wire_w_lg_read_sid_wire13w(0)) AND wire_w_lg_sec_protect_wire12w(0)) AND (NOT (read_wire OR fast_read_wire))) AND write_wire);
	do_write_polling <= wire_w_lg_w_lg_w661w806w807w(0);
	do_write_rstat <= write_rstat_reg;
	do_write_volatile <= '0';
	do_write_volatile_rstat <= '0';
	do_write_volatile_wren <= '0';
	do_write_wren <= ((NOT wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0));
	dummy_read_buf <= maxcnt_shift_reg2;
	end1_cyc_dlyncs_in_wire <= (((((((((wire_stage_cntr_w_lg_w_lg_w_q_range115w120w138w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND (NOT wire_gen_cntr_q(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range115w120w138w139w140w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w135w(0)) OR wire_w_lg_do_write84w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire130w(0)));
	end1_cyc_gen_cntr_wire <= (wire_gen_cntr_w_lg_w_q_range126w127w(0) AND (NOT wire_gen_cntr_q(0)));
	end1_cyc_normal_in_wire <= ((((((((((wire_stage_cntr_w_lg_w_lg_w_q_range115w120w138w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range115w120w138w139w140w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w135w(0)) OR wire_w_lg_do_write84w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire130w(0))) OR (do_read_rdid AND end_op_wire));
	end1_cyc_reg_in_wire <= wire_mux211_dataout;
	end_add_cycle <= wire_mux212_dataout;
	end_add_cycle_mux_datab_wire <= (wire_addbyte_cntr_q(2) AND wire_addbyte_cntr_q(1));
	end_fast_read <= end_read_reg;
	end_one_cyc_pos <= end1_cyc_reg2;
	end_one_cycle <= end1_cyc_reg;
	end_op_wire <= (((((((((((wire_stage_cntr_w_lg_w_q_range116w121w(0) AND ((wire_w_lg_w_lg_w_lg_w_lg_do_read394w395w396w397w(0) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read))) OR (wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w119w389w390w(0) AND wire_w_lg_do_polling219w(0))) OR ((((((do_read_rdid AND end_one_cyc_pos) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) AND wire_addbyte_cntr_q(2)) AND wire_addbyte_cntr_q(1)) AND wire_addbyte_cntr_w_lg_w_q_range177w178w(0))) OR (wire_w_lg_w_lg_start_poll380w381w(0) AND wire_w_lg_st_busy_wire130w(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range116w117w118w378w379w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write86w133w134w135w(0)) OR wire_w_lg_w_lg_do_write77w373w(0)) OR wire_w_lg_do_write84w(0)) OR wire_stage_cntr_w372w(0)) OR wire_stage_cntr_w_lg_w367w368w(0)) OR (wire_stage_cntr_w_lg_w_lg_w_q_range116w119w362w(0) AND ((do_write_volatile OR do_read_volatile) OR wire_w_lg_do_read_nonvolatile360w(0))));
	end_operation <= end_op_reg;
	end_ophdly <= end_op_hdlyreg;
	end_pgwr_data <= end_pgwrop_reg;
	end_read <= end_read_reg;
	end_read_byte <= (end_rbyte_reg AND wire_w_lg_addr_overdie539w(0));
	end_wrstage <= end_operation;
	exb4addr_opcode <= (OTHERS => '0');
	fast_read_opcode <= "00001011";
	fast_read_wire <= fast_read_reg;
	freadwrv_sdoin <= '0';
	ill_erase_wire <= ill_erase_reg;
	ill_write_wire <= ill_write_reg;
	illegal_erase <= ill_erase_wire;
	illegal_erase_b4out_wire <= (((do_sec_erase OR do_bulk_erase) OR do_die_erase) AND write_prot_true);
	illegal_write <= ill_write_wire;
	illegal_write_b4out_wire <= ((do_write AND write_prot_true) OR wire_w_lg_do_write84w(0));
	in_operation <= busy_wire;
	load_opcode <= ((((wire_stage_cntr_w_lg_w_q_range116w117w(0) AND wire_stage_cntr_w_lg_w_q_range115w120w(0)) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_w_lg_w_q_range124w125w(0)) AND wire_gen_cntr_q(0));
	mask_prot <= ( wire_w_lg_w707w709w & wire_w707w & wire_w_lg_w_lg_w_lg_w_prot_wire_range683w701w703w705w & wire_w_lg_w_lg_w_prot_wire_range683w701w703w & wire_w_lg_w_prot_wire_range683w701w & prot_wire(1));
	mask_prot_add <= ( wire_w_lg_w_mask_prot_range710w738w & wire_w_lg_w_mask_prot_range708w734w & wire_w_lg_w_mask_prot_range706w729w & wire_w_lg_w_mask_prot_range704w724w & wire_w_lg_w_mask_prot_range702w719w & wire_w_lg_w_mask_prot_range699w712w);
	mask_prot_check <= ( wire_w_lg_w_mask_prot_range710w740w & wire_w_lg_w_mask_prot_range708w736w & wire_w_lg_w_mask_prot_range706w731w & wire_w_lg_w_mask_prot_range704w726w & wire_w_lg_w_mask_prot_range702w721w & wire_w_lg_w_mask_prot_range699w715w);
	mask_prot_comp_ntb <= ( wire_w_lg_w_mask_prot_check_range741w762w & wire_w_lg_w_mask_prot_check_range737w758w & wire_w_lg_w_mask_prot_check_range732w754w & wire_w_lg_w_mask_prot_check_range727w750w & wire_w_lg_w_mask_prot_check_range722w746w & mask_prot_check(0));
	mask_prot_comp_tb <= ( wire_w_lg_w_mask_prot_add_range739w764w & wire_w_lg_w_mask_prot_add_range735w760w & wire_w_lg_w_mask_prot_add_range730w756w & wire_w_lg_w_mask_prot_add_range725w752w & wire_w_lg_w_mask_prot_add_range720w748w & mask_prot_add(0));
	memadd_sdoin <= add_msb_reg;
	ncs_reg_ena_wire <= (((wire_stage_cntr_w_lg_w_lg_w_q_range116w117w118w(0) AND end_one_cyc_pos) OR addr_overdie_pos) OR end_operation);
	not_busy <= busy_det_reg;
	oe_wire <= '0';
	page_size_wire <= "100000000";
	pagewr_buf_not_empty <= ( wire_w_lg_w_pagewr_buf_not_empty_range634w636w & wire_w_lg_w_pagewr_buf_not_empty_range631w633w & wire_w_lg_w_pagewr_buf_not_empty_range628w630w & wire_w_lg_w_pagewr_buf_not_empty_range625w627w & wire_w_lg_w_pagewr_buf_not_empty_range622w624w & wire_w_lg_w_pagewr_buf_not_empty_range619w621w & wire_w_lg_w_pagewr_buf_not_empty_range616w618w & wire_w_lg_w_pagewr_buf_not_empty_range612w615w & wire_pgwr_data_cntr_q(0));
	prot_wire <= ( wire_w_lg_w_lg_bp2_wire694w697w & wire_w_lg_w_lg_bp2_wire694w695w & wire_w_lg_w_lg_bp2_wire689w692w & wire_w_lg_w_lg_bp2_wire689w690w & wire_w_lg_w_lg_w_lg_bp2_wire677w684w687w & wire_w_lg_w_lg_w_lg_bp2_wire677w684w685w & wire_w_lg_w_lg_w_lg_bp2_wire677w678w682w & wire_w_lg_w_lg_w_lg_bp2_wire677w678w679w);
	rden_wire <= rden;
	rdid_load <= (end_operation AND do_read_rdid);
	rdid_opcode <= "10011111";
	rdid_out <= ( rdid_out_reg(7 DOWNTO 0));
	rdummyclk_opcode <= (OTHERS => '0');
	reach_max_cnt <= max_cnt_reg;
	read_address <= ( read_add_reg(23 DOWNTO 0));
	read_buf <= (((((end_one_cycle AND do_write) AND wire_w_lg_do_read_stat66w(0)) AND wire_w_lg_do_wren67w(0)) AND (wire_stage_cntr_w_lg_w_q_range116w121w(0) OR wire_addbyte_cntr_w_lg_w_q_range174w179w(0))) AND wire_w_lg_buf_empty780w(0));
	read_bufdly <= read_bufdly_reg;
	read_data_reg_in_wire <= ( read_dout_reg(7 DOWNTO 0));
	read_opcode <= (OTHERS => '0');
	read_rdid_wire <= read_rdid_reg;
	read_sid_wire <= '0';
	read_status_wire <= read_status_reg;
	read_wire <= '0';
	rflagstat_opcode <= "00000101";
	rnvdummyclk_opcode <= (OTHERS => '0');
	rsid_opcode <= (OTHERS => '0');
	rsid_sdoin <= '0';
	rstat_opcode <= "00000101";
	scein_wire <= wire_ncs_reg_w_lg_q415w(0);
	sdoin_wire <= to_sdoin_wire;
	sec_erase_wire <= sec_erase_reg;
	sec_protect_wire <= '0';
	secprot_opcode <= (OTHERS => '0');
	secprot_sdoin <= '0';
	serase_opcode <= "11011000";
	shift_bytes_wire <= shift_bytes;
	shift_opcode <= shift_op_reg;
	shift_opdata <= stage2_wire;
	shift_pgwr_data <= shftpgwr_data_reg;
	st_busy_wire <= statreg_int(0);
	stage2_wire <= stage2_reg;
	stage3_wire <= stage3_reg;
	stage4_wire <= stage4_reg;
	start_frpoll <= '0';
	start_poll <= ((start_wrpoll OR start_sppoll) OR start_frpoll);
	start_sppoll <= '0';
	start_wrpoll <= start_wrpoll_reg2;
	status_out <= ( statreg_out(7 DOWNTO 0));
	to_sdoin_wire <= ((((((shift_opdata AND asmi_opcode_reg(7)) OR rsid_sdoin) OR memadd_sdoin) OR write_sdoin) OR secprot_sdoin) OR freadwrv_sdoin);
	wren_opcode <= "00000110";
	wren_wire <= '1';
	write_opcode <= "00000010";
	write_prot_true <= write_prot_reg;
	write_sdoin <= ((((do_write AND stage4_wire) AND wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0)) AND pgwrbuf_dataout(7));
	write_wire <= write_reg;
	wrvolatile_opcode <= (OTHERS => '0');
	wire_w_addr_range438w(0) <= addr(0);
	wire_w_addr_range430w <= addr(23 DOWNTO 1);
	wire_w_addr_reg_overdie_range436w(0) <= addr_reg_overdie(0);
	wire_w_addr_reg_overdie_range426w <= addr_reg_overdie(23 DOWNTO 1);
	wire_w_b4addr_opcode_range282w(0) <= b4addr_opcode(0);
	wire_w_b4addr_opcode_range191w <= b4addr_opcode(7 DOWNTO 1);
	wire_w_berase_opcode_range286w(0) <= berase_opcode(0);
	wire_w_berase_opcode_range199w <= berase_opcode(7 DOWNTO 1);
	wire_w_dataout_wire_range478w(0) <= dataout_wire(1);
	wire_w_derase_opcode_range288w(0) <= derase_opcode(0);
	wire_w_derase_opcode_range204w <= derase_opcode(7 DOWNTO 1);
	wire_w_exb4addr_opcode_range280w(0) <= exb4addr_opcode(0);
	wire_w_exb4addr_opcode_range186w <= exb4addr_opcode(7 DOWNTO 1);
	wire_w_fast_read_opcode_range304w(0) <= fast_read_opcode(0);
	wire_w_fast_read_opcode_range244w <= fast_read_opcode(7 DOWNTO 1);
	wire_w_mask_prot_range699w(0) <= mask_prot(0);
	wire_w_mask_prot_range702w(0) <= mask_prot(1);
	wire_w_mask_prot_range704w(0) <= mask_prot(2);
	wire_w_mask_prot_range706w(0) <= mask_prot(3);
	wire_w_mask_prot_range708w(0) <= mask_prot(4);
	wire_w_mask_prot_range710w(0) <= mask_prot(5);
	wire_w_mask_prot_add_range713w(0) <= mask_prot_add(0);
	wire_w_mask_prot_add_range720w(0) <= mask_prot_add(1);
	wire_w_mask_prot_add_range725w(0) <= mask_prot_add(2);
	wire_w_mask_prot_add_range730w(0) <= mask_prot_add(3);
	wire_w_mask_prot_add_range735w(0) <= mask_prot_add(4);
	wire_w_mask_prot_add_range739w(0) <= mask_prot_add(5);
	wire_w_mask_prot_check_range722w(0) <= mask_prot_check(1);
	wire_w_mask_prot_check_range727w(0) <= mask_prot_check(2);
	wire_w_mask_prot_check_range732w(0) <= mask_prot_check(3);
	wire_w_mask_prot_check_range737w(0) <= mask_prot_check(4);
	wire_w_mask_prot_check_range741w(0) <= mask_prot_check(5);
	wire_w_mask_prot_comp_ntb_range742w(0) <= mask_prot_comp_ntb(0);
	wire_w_mask_prot_comp_ntb_range747w(0) <= mask_prot_comp_ntb(1);
	wire_w_mask_prot_comp_ntb_range751w(0) <= mask_prot_comp_ntb(2);
	wire_w_mask_prot_comp_ntb_range755w(0) <= mask_prot_comp_ntb(3);
	wire_w_mask_prot_comp_ntb_range759w(0) <= mask_prot_comp_ntb(4);
	wire_w_mask_prot_comp_tb_range744w(0) <= mask_prot_comp_tb(0);
	wire_w_mask_prot_comp_tb_range749w(0) <= mask_prot_comp_tb(1);
	wire_w_mask_prot_comp_tb_range753w(0) <= mask_prot_comp_tb(2);
	wire_w_mask_prot_comp_tb_range757w(0) <= mask_prot_comp_tb(3);
	wire_w_mask_prot_comp_tb_range761w(0) <= mask_prot_comp_tb(4);
	wire_w_pagewr_buf_not_empty_range612w(0) <= pagewr_buf_not_empty(0);
	wire_w_pagewr_buf_not_empty_range616w(0) <= pagewr_buf_not_empty(1);
	wire_w_pagewr_buf_not_empty_range619w(0) <= pagewr_buf_not_empty(2);
	wire_w_pagewr_buf_not_empty_range622w(0) <= pagewr_buf_not_empty(3);
	wire_w_pagewr_buf_not_empty_range625w(0) <= pagewr_buf_not_empty(4);
	wire_w_pagewr_buf_not_empty_range628w(0) <= pagewr_buf_not_empty(5);
	wire_w_pagewr_buf_not_empty_range631w(0) <= pagewr_buf_not_empty(6);
	wire_w_pagewr_buf_not_empty_range634w(0) <= pagewr_buf_not_empty(7);
	wire_w_pagewr_buf_not_empty_range82w(0) <= pagewr_buf_not_empty(8);
	wire_w_prot_wire_range683w(0) <= prot_wire(1);
	wire_w_prot_wire_range686w(0) <= prot_wire(2);
	wire_w_prot_wire_range688w(0) <= prot_wire(3);
	wire_w_prot_wire_range691w(0) <= prot_wire(4);
	wire_w_prot_wire_range693w(0) <= prot_wire(5);
	wire_w_prot_wire_range696w(0) <= prot_wire(6);
	wire_w_rdid_opcode_range310w(0) <= rdid_opcode(0);
	wire_w_rdid_opcode_range255w <= rdid_opcode(7 DOWNTO 1);
	wire_w_rdummyclk_opcode_range302w(0) <= rdummyclk_opcode(0);
	wire_w_rdummyclk_opcode_range237w <= rdummyclk_opcode(7 DOWNTO 1);
	wire_w_read_opcode_range306w(0) <= read_opcode(0);
	wire_w_read_opcode_range247w <= read_opcode(7 DOWNTO 1);
	wire_w_rflagstat_opcode_range292w(0) <= rflagstat_opcode(0);
	wire_w_rflagstat_opcode_range214w <= rflagstat_opcode(7 DOWNTO 1);
	wire_w_rnvdummyclk_opcode_range298w(0) <= rnvdummyclk_opcode(0);
	wire_w_rnvdummyclk_opcode_range227w <= rnvdummyclk_opcode(7 DOWNTO 1);
	wire_w_rsid_opcode_range312w(0) <= rsid_opcode(0);
	wire_w_rsid_opcode_range258w <= rsid_opcode(7 DOWNTO 1);
	wire_w_rstat_opcode_range294w(0) <= rstat_opcode(0);
	wire_w_rstat_opcode_range218w <= rstat_opcode(7 DOWNTO 1);
	wire_w_secprot_opcode_range308w(0) <= secprot_opcode(0);
	wire_w_secprot_opcode_range250w <= secprot_opcode(7 DOWNTO 1);
	wire_w_serase_opcode_range290w(0) <= serase_opcode(0);
	wire_w_serase_opcode_range209w <= serase_opcode(7 DOWNTO 1);
	wire_w_wren_opcode_range284w(0) <= wren_opcode(0);
	wire_w_wren_opcode_range196w <= wren_opcode(7 DOWNTO 1);
	wire_w_write_opcode_range296w(0) <= write_opcode(0);
	wire_w_write_opcode_range222w <= write_opcode(7 DOWNTO 1);
	wire_w_wrvolatile_opcode_range300w(0) <= wrvolatile_opcode(0);
	wire_w_wrvolatile_opcode_range230w <= wrvolatile_opcode(7 DOWNTO 1);
	wire_addbyte_cntr_w_lg_w_q_range174w179w(0) <= wire_addbyte_cntr_w_q_range174w(0) AND wire_addbyte_cntr_w_lg_w_q_range177w178w(0);
	wire_addbyte_cntr_w_lg_w_q_range177w178w(0) <= NOT wire_addbyte_cntr_w_q_range177w(0);
	wire_addbyte_cntr_clk_en <= wire_stage_cntr_w173w(0);
	wire_stage_cntr_w173w(0) <= ((wire_stage_cntr_w_lg_w_lg_w_q_range116w119w170w(0) AND wire_w_lg_w_lg_w167w168w169w(0)) OR addr_overdie) OR end_operation;
	wire_addbyte_cntr_clock <= wire_w_lg_clkin_wire48w(0);
	wire_addbyte_cntr_sclr <= wire_w_lg_end_operation114w(0);
	wire_w_lg_end_operation114w(0) <= end_operation OR addr_overdie;
	wire_addbyte_cntr_w_q_range177w(0) <= wire_addbyte_cntr_q(0);
	wire_addbyte_cntr_w_q_range174w(0) <= wire_addbyte_cntr_q(1);
	addbyte_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_addbyte_cntr_clk_en,
		clock => wire_addbyte_cntr_clock,
		q => wire_addbyte_cntr_q,
		sclr => wire_addbyte_cntr_sclr
	  );
	wire_gen_cntr_w_lg_w_q_range126w127w(0) <= wire_gen_cntr_w_q_range126w(0) AND wire_gen_cntr_w_lg_w_q_range124w125w(0);
	wire_gen_cntr_w_lg_w_q_range124w125w(0) <= NOT wire_gen_cntr_w_q_range124w(0);
	wire_gen_cntr_clk_en <= wire_w56w(0);
	wire_w56w(0) <= (((wire_w_lg_in_operation52w(0) AND wire_w_lg_clr_rstat_wire50w(0)) AND wire_w_lg_clr_sid_wire49w(0)) OR do_wait_dummyclk) OR addr_overdie;
	wire_gen_cntr_sclr <= wire_w_lg_w_lg_end1_cyc_reg_in_wire57w58w(0);
	wire_w_lg_w_lg_end1_cyc_reg_in_wire57w58w(0) <= (end1_cyc_reg_in_wire OR addr_overdie) OR do_wait_dummyclk;
	wire_gen_cntr_w_q_range124w(0) <= wire_gen_cntr_q(1);
	wire_gen_cntr_w_q_range126w(0) <= wire_gen_cntr_q(2);
	gen_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_gen_cntr_clk_en,
		clock => clkin_wire,
		q => wire_gen_cntr_q,
		sclr => wire_gen_cntr_sclr
	  );
	wire_stage_cntr_w_lg_w367w368w(0) <= wire_stage_cntr_w367w(0) AND end_one_cycle;
	wire_stage_cntr_w367w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range116w119w364w365w366w(0) AND end_add_cycle;
	wire_stage_cntr_w372w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range116w119w369w370w371w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range116w119w364w365w366w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w119w364w365w(0) AND wire_w_lg_do_read_stat66w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range116w119w369w370w371w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w119w369w370w(0) AND wire_w_lg_do_read_stat66w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range116w117w118w378w379w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w117w118w378w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w121w454w455w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range116w121w454w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w119w364w365w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range116w119w364w(0) AND wire_w_lg_do_wren67w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w119w389w390w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range116w119w389w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w119w369w370w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range116w119w369w(0) AND wire_w_lg_do_wren67w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range116w117w118w378w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range116w117w118w(0) AND wire_w_lg_do_wren377w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range116w121w454w(0) <= wire_stage_cntr_w_lg_w_q_range116w121w(0) AND end_add_cycle;
	wire_stage_cntr_w_lg_w_lg_w_q_range116w119w364w(0) <= wire_stage_cntr_w_lg_w_q_range116w119w(0) AND wire_w_lg_do_sec_erase68w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range116w119w389w(0) <= wire_stage_cntr_w_lg_w_q_range116w119w(0) AND do_read_stat;
	wire_stage_cntr_w_lg_w_lg_w_q_range116w119w369w(0) <= wire_stage_cntr_w_lg_w_q_range116w119w(0) AND do_sec_prot;
	wire_stage_cntr_w_lg_w_lg_w_q_range116w119w170w(0) <= wire_stage_cntr_w_lg_w_q_range116w119w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_q_range116w119w362w(0) <= wire_stage_cntr_w_lg_w_q_range116w119w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range115w120w138w139w140w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range115w120w138w139w(0) AND end1_cyc_gen_cntr_wire;
	wire_stage_cntr_w_lg_w_lg_w_q_range115w120w138w(0) <= wire_stage_cntr_w_lg_w_q_range115w120w(0) AND wire_stage_cntr_w_lg_w_q_range116w117w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range116w117w118w(0) <= wire_stage_cntr_w_lg_w_q_range116w117w(0) AND wire_stage_cntr_w_q_range115w(0);
	wire_stage_cntr_w_lg_w_q_range116w121w(0) <= wire_stage_cntr_w_q_range116w(0) AND wire_stage_cntr_w_lg_w_q_range115w120w(0);
	wire_stage_cntr_w_lg_w_q_range116w119w(0) <= wire_stage_cntr_w_q_range116w(0) AND wire_stage_cntr_w_q_range115w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range115w120w138w139w(0) <= NOT wire_stage_cntr_w_lg_w_lg_w_q_range115w120w138w(0);
	wire_stage_cntr_w_lg_w_q_range115w120w(0) <= NOT wire_stage_cntr_w_q_range115w(0);
	wire_stage_cntr_w_lg_w_q_range116w117w(0) <= NOT wire_stage_cntr_w_q_range116w(0);
	wire_stage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w110w111w112w113w(0);
	wire_w_lg_w_lg_w_lg_w110w111w112w113w(0) <= (((((((((((((in_operation AND end_one_cycle) AND (NOT (stage3_wire AND wire_w_lg_end_add_cycle97w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_read94w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_fast_read91w(0)))) AND (NOT ((wire_w_lg_w_lg_do_write86w87w(0) OR do_bulk_erase) AND write_prot_true))) AND (NOT wire_w_lg_do_write84w(0))) AND (NOT (stage3_wire AND st_busy_wire))) AND (NOT (wire_w_lg_do_write77w(0) AND wire_w_lg_end_pgwr_data76w(0)))) AND (NOT (stage2_wire AND do_wren))) AND (NOT (((wire_w_lg_stage3_wire69w(0) AND wire_w_lg_do_wren67w(0)) AND wire_w_lg_do_read_stat66w(0)) AND wire_w_lg_do_read_rdid65w(0)))) AND (NOT (stage3_wire AND ((do_write_volatile OR do_read_volatile) OR do_read_nonvolatile)))) OR wire_w_lg_w_lg_stage3_wire59w60w(0)) OR addr_overdie) OR end_ophdly;
	wire_stage_cntr_sclr <= wire_w_lg_end_operation114w(0);
	wire_stage_cntr_w_q_range115w(0) <= wire_stage_cntr_q(0);
	wire_stage_cntr_w_q_range116w(0) <= wire_stage_cntr_q(1);
	stage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_stage_cntr_clk_en,
		clock => clkin_wire,
		q => wire_stage_cntr_q,
		sclr => wire_stage_cntr_sclr
	  );
	wire_wrstage_cntr_w_lg_w_q_range655w656w(0) <= wire_wrstage_cntr_w_q_range655w(0) AND wire_wrstage_cntr_w_lg_w_q_range653w654w(0);
	wire_wrstage_cntr_w_lg_w_q_range653w654w(0) <= NOT wire_wrstage_cntr_w_q_range653w(0);
	wire_wrstage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w_lg_w648w649w650w651w652w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w648w649w650w651w652w(0) <= (wire_w_lg_w_lg_w648w649w650w(0) AND wire_w_lg_st_busy_wire130w(0)) OR clr_write_wire2;
	wire_wrstage_cntr_clock <= wire_w_lg_clkin_wire48w(0);
	wire_wrstage_cntr_w_q_range653w(0) <= wire_wrstage_cntr_q(0);
	wire_wrstage_cntr_w_q_range655w(0) <= wire_wrstage_cntr_q(1);
	wrstage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_wrstage_cntr_clk_en,
		clock => wire_wrstage_cntr_clock,
		q => wire_wrstage_cntr_q,
		sclr => clr_write_wire2
	  );
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN add_msb_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_add_msb_reg_ena = '1') THEN 
				IF (clr_addmsb_wire = '1') THEN add_msb_reg <= '0';
				ELSE add_msb_reg <= wire_addr_reg_w_q_range458w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_add_msb_reg_ena <= ((((wire_w_lg_w_lg_w_lg_w_lg_do_read335w462w463w464w(0) AND (NOT (wire_w_lg_w_lg_do_write86w87w(0) AND wire_w_lg_do_memadd459w(0)))) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) OR clr_addmsb_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN add_rollover_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN add_rollover_reg <= (wire_read_add_cntr_q(24) OR clr_read_wire2);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(0) = '1') THEN addr_reg(0) <= wire_addr_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(1) = '1') THEN addr_reg(1) <= wire_addr_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(2) = '1') THEN addr_reg(2) <= wire_addr_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(3) = '1') THEN addr_reg(3) <= wire_addr_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(4) = '1') THEN addr_reg(4) <= wire_addr_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(5) = '1') THEN addr_reg(5) <= wire_addr_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(6) = '1') THEN addr_reg(6) <= wire_addr_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(7) = '1') THEN addr_reg(7) <= wire_addr_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(8) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(8) = '1') THEN addr_reg(8) <= wire_addr_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(9) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(9) = '1') THEN addr_reg(9) <= wire_addr_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(10) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(10) = '1') THEN addr_reg(10) <= wire_addr_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(11) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(11) = '1') THEN addr_reg(11) <= wire_addr_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(12) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(12) = '1') THEN addr_reg(12) <= wire_addr_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(13) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(13) = '1') THEN addr_reg(13) <= wire_addr_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(14) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(14) = '1') THEN addr_reg(14) <= wire_addr_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(15) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(15) = '1') THEN addr_reg(15) <= wire_addr_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(16) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(16) = '1') THEN addr_reg(16) <= wire_addr_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(17) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(17) = '1') THEN addr_reg(17) <= wire_addr_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(18) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(18) = '1') THEN addr_reg(18) <= wire_addr_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(19) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(19) = '1') THEN addr_reg(19) <= wire_addr_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(20) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(20) = '1') THEN addr_reg(20) <= wire_addr_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(21) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(21) = '1') THEN addr_reg(21) <= wire_addr_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(22) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(22) = '1') THEN addr_reg(22) <= wire_addr_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(23) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(23) = '1') THEN addr_reg(23) <= wire_addr_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_addr_reg_d <= ( wire_w_lg_w_lg_w_lg_not_busy431w432w433w & wire_w_lg_w_lg_not_busy439w440w);
	loop43 : FOR i IN 0 TO 23 GENERATE
		wire_addr_reg_ena(i) <= wire_w_lg_w_lg_w_lg_w_lg_rden_wire446w447w448w449w(0);
	END GENERATE loop43;
	wire_addr_reg_w_q_range711w(0) <= addr_reg(18);
	wire_addr_reg_w_q_range718w(0) <= addr_reg(19);
	wire_addr_reg_w_q_range723w(0) <= addr_reg(20);
	wire_addr_reg_w_q_range728w(0) <= addr_reg(21);
	wire_addr_reg_w_q_range428w <= addr_reg(22 DOWNTO 0);
	wire_addr_reg_w_q_range733w(0) <= addr_reg(22);
	wire_addr_reg_w_q_range458w(0) <= addr_reg(23);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(0) = '1') THEN asmi_opcode_reg(0) <= wire_asmi_opcode_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(1) = '1') THEN asmi_opcode_reg(1) <= wire_asmi_opcode_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(2) = '1') THEN asmi_opcode_reg(2) <= wire_asmi_opcode_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(3) = '1') THEN asmi_opcode_reg(3) <= wire_asmi_opcode_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(4) = '1') THEN asmi_opcode_reg(4) <= wire_asmi_opcode_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(5) = '1') THEN asmi_opcode_reg(5) <= wire_asmi_opcode_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(6) = '1') THEN asmi_opcode_reg(6) <= wire_asmi_opcode_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(7) = '1') THEN asmi_opcode_reg(7) <= wire_asmi_opcode_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_asmi_opcode_reg_d <= ( wire_w_lg_w_lg_w275w276w277w & wire_w_lg_w328w329w);
	loop44 : FOR i IN 0 TO 7 GENERATE
		wire_asmi_opcode_reg_ena(i) <= wire_w_lg_load_opcode331w(0);
	END GENERATE loop44;
	wire_asmi_opcode_reg_w_q_range184w <= asmi_opcode_reg(6 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN buf_empty_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN buf_empty_reg <= wire_cmpr5_aeb;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN busy_delay_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (power_up_reg = '1') THEN busy_delay_reg <= busy_wire;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN busy_det_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN busy_det_reg <= wire_w_lg_busy_wire3w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_rdid_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rdid_reg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_read_reg <= ((do_read_sid OR do_sec_prot) OR wire_w_lg_end_operation545w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN clr_read_reg2 <= clr_read_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_rstat_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN clr_rstat_reg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_write_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_write_reg <= ((((((wire_w_lg_w_lg_w_lg_w_lg_w661w806w807w817w818w(0) OR wire_w_lg_do_write84w(0)) OR wire_w_lg_w_lg_w814w815w816w(0)) OR do_read_sid) OR do_sec_prot) OR do_read) OR do_fast_read);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_write_reg2 <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_write_reg2 <= clr_write_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN cnt_bfend_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN cnt_bfend_reg <= cnt_bfend_wire_in;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN do_wrmemadd_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN do_wrmemadd_reg <= (wire_wrstage_cntr_q(1) AND wire_wrstage_cntr_q(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_dvalid_reg_ena = '1') THEN 
				IF (wire_dvalid_reg_sclr = '1') THEN dvalid_reg <= '0';
				ELSE dvalid_reg <= wire_w_lg_end_read_byte514w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_dvalid_reg_ena <= wire_w_lg_do_read335w(0);
	wire_dvalid_reg_sclr <= (end_op_wire OR end_operation);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN dvalid_reg2 <= dvalid_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end1_cyc_reg <= end1_cyc_reg_in_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end1_cyc_reg2 <= end_one_cycle;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_hdlyreg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_op_hdlyreg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end_op_reg <= end_op_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_pgwrop_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_end_pgwrop_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN end_pgwrop_reg <= '0';
				ELSE end_pgwrop_reg <= buf_empty;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_end_pgwrop_reg_ena <= (((cnt_bfend_reg AND do_write) AND shift_pgwr_data) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_rbyte_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_end_rbyte_reg_ena = '1') THEN 
				IF (wire_end_rbyte_reg_sclr = '1') THEN end_rbyte_reg <= '0';
				ELSE end_rbyte_reg <= wire_w_lg_w_lg_w_lg_do_read335w507w508w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_end_rbyte_reg_ena <= ((wire_gen_cntr_w_lg_w_q_range126w127w(0) AND wire_gen_cntr_q(0)) OR clr_endrbyte_wire);
	wire_end_rbyte_reg_sclr <= (clr_endrbyte_wire OR addr_overdie);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_read_reg <= (((wire_w_lg_rden_wire541w(0) AND wire_w_lg_do_read335w(0)) AND data_valid_wire) AND end_read_byte);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN fast_read_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_fast_read_reg_ena = '1') THEN 
				IF (clr_read_wire = '1') THEN fast_read_reg <= '0';
				ELSE fast_read_reg <= fast_read;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_fast_read_reg_ena <= ((wire_w_lg_busy_wire3w(0) AND rden_wire) OR clr_read_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN ill_erase_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN ill_erase_reg <= (illegal_erase_dly_reg OR illegal_erase_b4out_wire);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN ill_write_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN ill_write_reg <= (illegal_write_dly_reg OR illegal_write_b4out_wire);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN illegal_erase_dly_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (power_up_reg = '1') THEN illegal_erase_dly_reg <= illegal_erase_b4out_wire;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN illegal_write_dly_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (power_up_reg = '1') THEN illegal_write_dly_reg <= illegal_write_b4out_wire;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN illegal_write_prot_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN illegal_write_prot_reg <= do_write;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN max_cnt_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN max_cnt_reg <= wire_cmpr4_aeb;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN maxcnt_shift_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN maxcnt_shift_reg <= (wire_w_lg_w_lg_reach_max_cnt643w644w(0) AND wire_w_lg_do_write563w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN maxcnt_shift_reg2 <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN maxcnt_shift_reg2 <= maxcnt_shift_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN ncs_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (ncs_reg_ena_wire = '1') THEN 
				IF (wire_ncs_reg_sclr = '1') THEN ncs_reg <= '0';
				ELSE ncs_reg <= '1';
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_ncs_reg_sclr <= (end_operation OR addr_overdie_pos);
	wire_ncs_reg_w_lg_q415w(0) <= NOT ncs_reg;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(0) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(0) <= '0';
				ELSE pgwrbuf_dataout(0) <= wire_pgwrbuf_dataout_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(1) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(1) <= '0';
				ELSE pgwrbuf_dataout(1) <= wire_pgwrbuf_dataout_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(2) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(2) <= '0';
				ELSE pgwrbuf_dataout(2) <= wire_pgwrbuf_dataout_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(3) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(3) <= '0';
				ELSE pgwrbuf_dataout(3) <= wire_pgwrbuf_dataout_d(3);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(4) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(4) <= '0';
				ELSE pgwrbuf_dataout(4) <= wire_pgwrbuf_dataout_d(4);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(5) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(5) <= '0';
				ELSE pgwrbuf_dataout(5) <= wire_pgwrbuf_dataout_d(5);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(6) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(6) <= '0';
				ELSE pgwrbuf_dataout(6) <= wire_pgwrbuf_dataout_d(6);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(7) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(7) <= '0';
				ELSE pgwrbuf_dataout(7) <= wire_pgwrbuf_dataout_d(7);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_pgwrbuf_dataout_d <= ( wire_w_lg_w_lg_read_bufdly600w601w & wire_w_lg_read_bufdly605w);
	loop45 : FOR i IN 0 TO 7 GENERATE
		wire_pgwrbuf_dataout_ena(i) <= wire_w_lg_w_lg_read_bufdly594w595w(0);
	END GENERATE loop45;
	wire_pgwrbuf_dataout_w_q_range596w <= pgwrbuf_dataout(6 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN power_up_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN power_up_reg <= (busy_wire OR busy_delay_reg);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN rdid_out_reg <= (OTHERS => '0');
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (rdid_load = '1') THEN rdid_out_reg <= ( read_dout_reg(7 DOWNTO 0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(0) = '1') THEN read_add_reg(0) <= wire_read_add_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(1) = '1') THEN read_add_reg(1) <= wire_read_add_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(2) = '1') THEN read_add_reg(2) <= wire_read_add_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(3) = '1') THEN read_add_reg(3) <= wire_read_add_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(4) = '1') THEN read_add_reg(4) <= wire_read_add_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(5) = '1') THEN read_add_reg(5) <= wire_read_add_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(6) = '1') THEN read_add_reg(6) <= wire_read_add_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(7) = '1') THEN read_add_reg(7) <= wire_read_add_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(8) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(8) = '1') THEN read_add_reg(8) <= wire_read_add_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(9) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(9) = '1') THEN read_add_reg(9) <= wire_read_add_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(10) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(10) = '1') THEN read_add_reg(10) <= wire_read_add_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(11) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(11) = '1') THEN read_add_reg(11) <= wire_read_add_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(12) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(12) = '1') THEN read_add_reg(12) <= wire_read_add_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(13) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(13) = '1') THEN read_add_reg(13) <= wire_read_add_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(14) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(14) = '1') THEN read_add_reg(14) <= wire_read_add_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(15) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(15) = '1') THEN read_add_reg(15) <= wire_read_add_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(16) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(16) = '1') THEN read_add_reg(16) <= wire_read_add_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(17) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(17) = '1') THEN read_add_reg(17) <= wire_read_add_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(18) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(18) = '1') THEN read_add_reg(18) <= wire_read_add_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(19) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(19) = '1') THEN read_add_reg(19) <= wire_read_add_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(20) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(20) = '1') THEN read_add_reg(20) <= wire_read_add_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(21) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(21) = '1') THEN read_add_reg(21) <= wire_read_add_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(22) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(22) = '1') THEN read_add_reg(22) <= wire_read_add_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(23) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(23) = '1') THEN read_add_reg(23) <= wire_read_add_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_read_add_reg_d <= ( wire_read_add_cntr_q(23 DOWNTO 0));
	loop46 : FOR i IN 0 TO 23 GENERATE
		wire_read_add_reg_ena(i) <= wire_w_lg_w_lg_end_read_byte514w526w(0);
	END GENERATE loop46;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_bufdly_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN read_bufdly_reg <= read_buf;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(0) = '1') THEN read_data_reg(0) <= wire_read_data_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(1) = '1') THEN read_data_reg(1) <= wire_read_data_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(2) = '1') THEN read_data_reg(2) <= wire_read_data_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(3) = '1') THEN read_data_reg(3) <= wire_read_data_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(4) = '1') THEN read_data_reg(4) <= wire_read_data_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(5) = '1') THEN read_data_reg(5) <= wire_read_data_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(6) = '1') THEN read_data_reg(6) <= wire_read_data_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(7) = '1') THEN read_data_reg(7) <= wire_read_data_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_data_reg_d <= ( read_data_reg_in_wire(7 DOWNTO 0));
	loop47 : FOR i IN 0 TO 7 GENERATE
		wire_read_data_reg_ena(i) <= wire_w510w(0);
	END GENERATE loop47;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(0) = '1') THEN read_dout_reg(0) <= wire_read_dout_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(1) = '1') THEN read_dout_reg(1) <= wire_read_dout_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(2) = '1') THEN read_dout_reg(2) <= wire_read_dout_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(3) = '1') THEN read_dout_reg(3) <= wire_read_dout_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(4) = '1') THEN read_dout_reg(4) <= wire_read_dout_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(5) = '1') THEN read_dout_reg(5) <= wire_read_dout_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(6) = '1') THEN read_dout_reg(6) <= wire_read_dout_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(7) = '1') THEN read_dout_reg(7) <= wire_read_dout_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_dout_reg_d <= ( read_dout_reg(6 DOWNTO 0) & wire_w_lg_data0out_wire479w);
	loop48 : FOR i IN 0 TO 7 GENERATE
		wire_read_dout_reg_ena(i) <= wire_w_lg_w_lg_stage4_wire476w477w(0);
	END GENERATE loop48;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_rdid_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_rdid_reg_ena = '1') THEN 
				IF (clr_rdid_wire = '1') THEN read_rdid_reg <= '0';
				ELSE read_rdid_reg <= read_rdid;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_read_rdid_reg_ena <= (wire_w_lg_busy_wire3w(0) OR clr_rdid_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_status_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_status_reg_ena = '1') THEN 
				IF (clr_rstat_wire = '1') THEN read_status_reg <= '0';
				ELSE read_status_reg <= read_status;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_read_status_reg_ena <= (wire_w_lg_busy_wire3w(0) OR clr_rstat_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN sec_erase_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_sec_erase_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN sec_erase_reg <= '0';
				ELSE sec_erase_reg <= sector_erase;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_sec_erase_reg_ena <= ((wire_w_lg_busy_wire3w(0) AND wren_wire) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN shftpgwr_data_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
				IF (end_operation = '1') THEN shftpgwr_data_reg <= '0';
				ELSE shftpgwr_data_reg <= ((wire_stage_cntr_w_lg_w_q_range116w121w(0) AND wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0));
				END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN shift_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN shift_op_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range116w117w118w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage2_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage2_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range116w117w118w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage3_dly_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN stage3_dly_reg <= wire_stage_cntr_w_lg_w_q_range116w119w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage3_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage3_reg <= wire_stage_cntr_w_lg_w_q_range116w119w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage4_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage4_reg <= wire_stage_cntr_w_lg_w_q_range116w121w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN start_wrpoll_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_start_wrpoll_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN start_wrpoll_reg <= '0';
				ELSE start_wrpoll_reg <= wire_stage_cntr_w_lg_w_q_range116w119w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_start_wrpoll_reg_ena <= (((do_write_rstat AND do_polling) AND end_one_cycle) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN start_wrpoll_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
				IF (clr_write_wire = '1') THEN start_wrpoll_reg2 <= '0';
				ELSE start_wrpoll_reg2 <= start_wrpoll_reg;
				END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(0) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(0) <= '0';
				ELSE statreg_int(0) <= wire_statreg_int_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(1) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(1) <= '0';
				ELSE statreg_int(1) <= wire_statreg_int_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(2) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(2) <= '0';
				ELSE statreg_int(2) <= wire_statreg_int_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(3) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(3) <= '0';
				ELSE statreg_int(3) <= wire_statreg_int_d(3);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(4) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(4) <= '0';
				ELSE statreg_int(4) <= wire_statreg_int_d(4);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(5) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(5) <= '0';
				ELSE statreg_int(5) <= wire_statreg_int_d(5);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(6) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(6) <= '0';
				ELSE statreg_int(6) <= wire_statreg_int_d(6);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(7) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(7) <= '0';
				ELSE statreg_int(7) <= wire_statreg_int_d(7);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_statreg_int_d <= ( read_dout_reg(7 DOWNTO 0));
	loop49 : FOR i IN 0 TO 7 GENERATE
		wire_statreg_int_ena(i) <= wire_w_lg_w_lg_w_lg_end_operation579w580w581w(0);
	END GENERATE loop49;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(0) = '1') THEN statreg_out(0) <= wire_statreg_out_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(1) = '1') THEN statreg_out(1) <= wire_statreg_out_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(2) = '1') THEN statreg_out(2) <= wire_statreg_out_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(3) = '1') THEN statreg_out(3) <= wire_statreg_out_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(4) = '1') THEN statreg_out(4) <= wire_statreg_out_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(5) = '1') THEN statreg_out(5) <= wire_statreg_out_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(6) = '1') THEN statreg_out(6) <= wire_statreg_out_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(7) = '1') THEN statreg_out(7) <= wire_statreg_out_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_statreg_out_d <= ( read_dout_reg(7 DOWNTO 0));
	loop50 : FOR i IN 0 TO 7 GENERATE
		wire_statreg_out_ena(i) <= wire_w_lg_w_lg_w_lg_w568w569w570w571w(0);
	END GENERATE loop50;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN write_prot_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_write_prot_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN write_prot_reg <= '0';
				ELSE write_prot_reg <= (((wire_w_lg_do_write86w(0) AND (NOT mask_prot_comp_ntb(5))) AND (NOT prot_wire(0))) OR be_write_prot);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_write_prot_reg_ena <= ((((wire_w_lg_w_lg_w_lg_do_sec_erase663w664w665w(0) AND (NOT wire_wrstage_cntr_q(1))) AND wire_wrstage_cntr_q(0)) AND end_ophdly) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN write_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_write_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN write_reg <= '0';
				ELSE write_reg <= write;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_write_reg_ena <= ((wire_w_lg_busy_wire3w(0) AND wren_wire) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN write_rstat_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
				IF (clr_write_wire = '1') THEN write_rstat_reg <= '0';
				ELSE write_rstat_reg <= (wire_w661w(0) AND (((NOT wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_w_lg_w_q_range653w654w(0)) OR wire_wrstage_cntr_w_lg_w_q_range655w656w(0)));
				END IF;
		END IF;
	END PROCESS;
	wire_cmpr4_dataa <= ( page_size_wire(8 DOWNTO 0));
	wire_cmpr4_datab <= ( wire_pgwr_data_cntr_q(8 DOWNTO 0));
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aeb => wire_cmpr4_aeb,
		dataa => wire_cmpr4_dataa,
		datab => wire_cmpr4_datab
	  );
	wire_cmpr5_dataa <= ( wire_pgwr_data_cntr_q(8 DOWNTO 0));
	wire_cmpr5_datab <= ( wire_pgwr_read_cntr_q(8 DOWNTO 0));
	cmpr5 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aeb => wire_cmpr5_aeb,
		dataa => wire_cmpr5_dataa,
		datab => wire_cmpr5_datab
	  );
	wire_pgwr_data_cntr_clk_en <= wire_w610w(0);
	wire_w610w(0) <= (((shift_bytes_wire AND wren_wire) AND wire_w_lg_reach_max_cnt607w(0)) AND wire_w_lg_do_write563w(0)) OR clr_write_wire2;
	wire_pgwr_data_cntr_w_q_range614w(0) <= wire_pgwr_data_cntr_q(1);
	wire_pgwr_data_cntr_w_q_range617w(0) <= wire_pgwr_data_cntr_q(2);
	wire_pgwr_data_cntr_w_q_range620w(0) <= wire_pgwr_data_cntr_q(3);
	wire_pgwr_data_cntr_w_q_range623w(0) <= wire_pgwr_data_cntr_q(4);
	wire_pgwr_data_cntr_w_q_range626w(0) <= wire_pgwr_data_cntr_q(5);
	wire_pgwr_data_cntr_w_q_range629w(0) <= wire_pgwr_data_cntr_q(6);
	wire_pgwr_data_cntr_w_q_range632w(0) <= wire_pgwr_data_cntr_q(7);
	wire_pgwr_data_cntr_w_q_range635w(0) <= wire_pgwr_data_cntr_q(8);
	pgwr_data_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 9
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_pgwr_data_cntr_clk_en,
		clock => clkin_wire,
		q => wire_pgwr_data_cntr_q,
		sclr => clr_write_wire2
	  );
	wire_pgwr_read_cntr_clk_en <= wire_w_lg_read_buf789w(0);
	wire_w_lg_read_buf789w(0) <= read_buf OR clr_write_wire2;
	pgwr_read_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 9
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_pgwr_read_cntr_clk_en,
		clock => clkin_wire,
		q => wire_pgwr_read_cntr_q,
		sclr => clr_write_wire2
	  );
	wire_read_add_cntr_clk_en <= wire_w_lg_w_lg_w_lg_rden_wire516w517w518w(0);
	wire_w_lg_w_lg_w_lg_rden_wire516w517w518w(0) <= ((rden_wire AND not_busy) OR data_valid_wire) OR add_rollover;
	wire_read_add_cntr_data <= ( "0" & addr(23 DOWNTO 0));
	wire_read_add_cntr_sload <= wire_w_lg_rden_wire516w(0);
	wire_w_lg_rden_wire516w(0) <= rden_wire AND not_busy;
	read_add_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 25
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_read_add_cntr_clk_en,
		clock => clkin_wire,
		data => wire_read_add_cntr_data,
		q => wire_read_add_cntr_q,
		sclr => add_rollover,
		sload => wire_read_add_cntr_sload
	  );
	wire_mux211_dataout <= end1_cyc_dlyncs_in_wire WHEN ((((do_write OR do_sec_prot) OR do_sec_erase) OR do_bulk_erase) OR do_die_erase) = '1'  ELSE end1_cyc_normal_in_wire;
	wire_mux212_dataout <= end_add_cycle_mux_datab_wire WHEN do_fast_read = '1'  ELSE wire_addbyte_cntr_w_lg_w_q_range174w179w(0);
	wire_scfifo3_data <= ( datain(7 DOWNTO 0));
	wire_scfifo3_rdreq <= wire_w_lg_read_buf593w(0);
	wire_w_lg_read_buf593w(0) <= read_buf OR dummy_read_buf;
	wire_scfifo3_wrreq <= wire_w_lg_w_lg_shift_bytes_wire591w592w(0);
	wire_w_lg_w_lg_shift_bytes_wire591w592w(0) <= (shift_bytes_wire AND wren_wire) AND wire_w_lg_do_write563w(0);
	wire_scfifo3_w_q_range599w <= wire_scfifo3_q(7 DOWNTO 1);
	wire_scfifo3_w_q_range604w(0) <= wire_scfifo3_q(0);
	scfifo3 :  scfifo
	  GENERIC MAP (
		LPM_NUMWORDS => 258,
		LPM_WIDTH => 8,
		LPM_WIDTHU => 9,
		USE_EAB => "ON"
	  )
	  PORT MAP ( 
		aclr => reset,
		clock => clkin_wire,
		data => wire_scfifo3_data,
		q => wire_scfifo3_q,
		rdreq => wire_scfifo3_rdreq,
		sclr => clr_write_wire2,
		wrreq => wire_scfifo3_wrreq
	  );

 END RTL; --altasmi_altasmi_parallel_di43
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altasmi IS
	PORT
	(
		addr		: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		asmi_dataout		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		clkin		: IN STD_LOGIC ;
		datain		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		fast_read		: IN STD_LOGIC ;
		rden		: IN STD_LOGIC ;
		read_rdid		: IN STD_LOGIC ;
		read_status		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		sector_erase		: IN STD_LOGIC ;
		shift_bytes		: IN STD_LOGIC ;
		write		: IN STD_LOGIC ;
		asmi_dataoe		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		asmi_dclk		: OUT STD_LOGIC ;
		asmi_scein		: OUT STD_LOGIC ;
		asmi_sdoin		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		busy		: OUT STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		illegal_erase		: OUT STD_LOGIC ;
		illegal_write		: OUT STD_LOGIC ;
		rdid_out		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		read_address		: OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
		status_out		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END altasmi;


ARCHITECTURE RTL OF altasmi IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "ALTASMI_PARALLEL";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "data_width=STANDARD;enable_sim=FALSE;epcs_type=EPCS128;flash_rstpin=FALSE;intended_device_family=Arria II GX;lpm_hint=UNUSED;lpm_type=altasmi_parallel;page_size=256;port_bulk_erase=PORT_UNUSED;port_die_erase=PORT_UNUSED;port_en4b_addr=PORT_UNUSED;port_ex4b_addr=PORT_UNUSED;port_fast_read=PORT_USED;port_illegal_erase=PORT_USED;port_illegal_write=PORT_USED;port_rdid_out=PORT_USED;port_read_address=PORT_USED;port_read_dummyclk=PORT_UNUSED;port_read_rdid=PORT_USED;port_read_sid=PORT_UNUSED;port_read_status=PORT_USED;port_sector_erase=PORT_USED;port_sector_protect=PORT_UNUSED;port_shift_bytes=PORT_USED;port_wren=PORT_UNUSED;port_write=PORT_USED;use_asmiblock=OFF;use_eab=ON;write_dummy_clk=0;";
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC ;
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC ;
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC ;
	SIGNAL sub_wire8	: STD_LOGIC ;
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (23 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (7 DOWNTO 0);



	COMPONENT altasmi_altasmi_parallel_di43
	PORT (
			addr	: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
			asmi_dataout	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			clkin	: IN STD_LOGIC ;
			datain	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			fast_read	: IN STD_LOGIC ;
			rden	: IN STD_LOGIC ;
			read_rdid	: IN STD_LOGIC ;
			read_status	: IN STD_LOGIC ;
			reset	: IN STD_LOGIC ;
			sector_erase	: IN STD_LOGIC ;
			shift_bytes	: IN STD_LOGIC ;
			write	: IN STD_LOGIC ;
			asmi_dataoe	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			asmi_dclk	: OUT STD_LOGIC ;
			asmi_scein	: OUT STD_LOGIC ;
			asmi_sdoin	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			data_valid	: OUT STD_LOGIC ;
			dataout	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			illegal_erase	: OUT STD_LOGIC ;
			illegal_write	: OUT STD_LOGIC ;
			rdid_out	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			read_address	: OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
			status_out	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	asmi_dataoe    <= sub_wire0(0 DOWNTO 0);
	asmi_dclk    <= sub_wire1;
	asmi_scein    <= sub_wire2;
	asmi_sdoin    <= sub_wire3(0 DOWNTO 0);
	busy    <= sub_wire4;
	data_valid    <= sub_wire5;
	dataout    <= sub_wire6(7 DOWNTO 0);
	illegal_erase    <= sub_wire7;
	illegal_write    <= sub_wire8;
	rdid_out    <= sub_wire9(7 DOWNTO 0);
	read_address    <= sub_wire10(23 DOWNTO 0);
	status_out    <= sub_wire11(7 DOWNTO 0);

	altasmi_altasmi_parallel_di43_component : altasmi_altasmi_parallel_di43
	PORT MAP (
		addr => addr,
		asmi_dataout => asmi_dataout,
		clkin => clkin,
		datain => datain,
		fast_read => fast_read,
		rden => rden,
		read_rdid => read_rdid,
		read_status => read_status,
		reset => reset,
		sector_erase => sector_erase,
		shift_bytes => shift_bytes,
		write => write,
		asmi_dataoe => sub_wire0,
		asmi_dclk => sub_wire1,
		asmi_scein => sub_wire2,
		asmi_sdoin => sub_wire3,
		busy => sub_wire4,
		data_valid => sub_wire5,
		dataout => sub_wire6,
		illegal_erase => sub_wire7,
		illegal_write => sub_wire8,
		rdid_out => sub_wire9,
		read_address => sub_wire10,
		status_out => sub_wire11
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: CONSTANT: DATA_WIDTH STRING "STANDARD"
-- Retrieval info: CONSTANT: ENABLE_SIM STRING "FALSE"
-- Retrieval info: CONSTANT: EPCS_TYPE STRING "EPCS128"
-- Retrieval info: CONSTANT: FLASH_RSTPIN STRING "FALSE"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altasmi_parallel"
-- Retrieval info: CONSTANT: PAGE_SIZE NUMERIC "256"
-- Retrieval info: CONSTANT: PORT_BULK_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_DIE_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_EN4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_EX4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_FAST_READ STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_ERASE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_WRITE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_RDID_OUT STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_ADDRESS STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_DUMMYCLK STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_RDID STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_SID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_STATUS STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_SECTOR_ERASE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_SECTOR_PROTECT STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SHIFT_BYTES STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_WREN STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_WRITE STRING "PORT_USED"
-- Retrieval info: CONSTANT: USE_ASMIBLOCK STRING "OFF"
-- Retrieval info: CONSTANT: USE_EAB STRING "ON"
-- Retrieval info: CONSTANT: WRITE_DUMMY_CLK NUMERIC "0"
-- Retrieval info: USED_PORT: addr 0 0 24 0 INPUT NODEFVAL "addr[23..0]"
-- Retrieval info: CONNECT: @addr 0 0 24 0 addr 0 0 24 0
-- Retrieval info: USED_PORT: asmi_dataoe 0 0 1 0 OUTPUT NODEFVAL "asmi_dataoe[0..0]"
-- Retrieval info: CONNECT: asmi_dataoe 0 0 1 0 @asmi_dataoe 0 0 1 0
-- Retrieval info: USED_PORT: asmi_dataout 0 0 1 0 INPUT NODEFVAL "asmi_dataout[0..0]"
-- Retrieval info: CONNECT: @asmi_dataout 0 0 1 0 asmi_dataout 0 0 1 0
-- Retrieval info: USED_PORT: asmi_dclk 0 0 0 0 OUTPUT NODEFVAL "asmi_dclk"
-- Retrieval info: CONNECT: asmi_dclk 0 0 0 0 @asmi_dclk 0 0 0 0
-- Retrieval info: USED_PORT: asmi_scein 0 0 0 0 OUTPUT NODEFVAL "asmi_scein"
-- Retrieval info: CONNECT: asmi_scein 0 0 0 0 @asmi_scein 0 0 0 0
-- Retrieval info: USED_PORT: asmi_sdoin 0 0 1 0 OUTPUT NODEFVAL "asmi_sdoin[0..0]"
-- Retrieval info: CONNECT: asmi_sdoin 0 0 1 0 @asmi_sdoin 0 0 1 0
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: USED_PORT: clkin 0 0 0 0 INPUT NODEFVAL "clkin"
-- Retrieval info: CONNECT: @clkin 0 0 0 0 clkin 0 0 0 0
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: USED_PORT: datain 0 0 8 0 INPUT NODEFVAL "datain[7..0]"
-- Retrieval info: CONNECT: @datain 0 0 8 0 datain 0 0 8 0
-- Retrieval info: USED_PORT: dataout 0 0 8 0 OUTPUT NODEFVAL "dataout[7..0]"
-- Retrieval info: CONNECT: dataout 0 0 8 0 @dataout 0 0 8 0
-- Retrieval info: USED_PORT: fast_read 0 0 0 0 INPUT NODEFVAL "fast_read"
-- Retrieval info: CONNECT: @fast_read 0 0 0 0 fast_read 0 0 0 0
-- Retrieval info: USED_PORT: illegal_erase 0 0 0 0 OUTPUT NODEFVAL "illegal_erase"
-- Retrieval info: CONNECT: illegal_erase 0 0 0 0 @illegal_erase 0 0 0 0
-- Retrieval info: USED_PORT: illegal_write 0 0 0 0 OUTPUT NODEFVAL "illegal_write"
-- Retrieval info: CONNECT: illegal_write 0 0 0 0 @illegal_write 0 0 0 0
-- Retrieval info: USED_PORT: rden 0 0 0 0 INPUT NODEFVAL "rden"
-- Retrieval info: CONNECT: @rden 0 0 0 0 rden 0 0 0 0
-- Retrieval info: USED_PORT: rdid_out 0 0 8 0 OUTPUT NODEFVAL "rdid_out[7..0]"
-- Retrieval info: CONNECT: rdid_out 0 0 8 0 @rdid_out 0 0 8 0
-- Retrieval info: USED_PORT: read_address 0 0 24 0 OUTPUT NODEFVAL "read_address[23..0]"
-- Retrieval info: CONNECT: read_address 0 0 24 0 @read_address 0 0 24 0
-- Retrieval info: USED_PORT: read_rdid 0 0 0 0 INPUT NODEFVAL "read_rdid"
-- Retrieval info: CONNECT: @read_rdid 0 0 0 0 read_rdid 0 0 0 0
-- Retrieval info: USED_PORT: read_status 0 0 0 0 INPUT NODEFVAL "read_status"
-- Retrieval info: CONNECT: @read_status 0 0 0 0 read_status 0 0 0 0
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: USED_PORT: sector_erase 0 0 0 0 INPUT NODEFVAL "sector_erase"
-- Retrieval info: CONNECT: @sector_erase 0 0 0 0 sector_erase 0 0 0 0
-- Retrieval info: USED_PORT: shift_bytes 0 0 0 0 INPUT NODEFVAL "shift_bytes"
-- Retrieval info: CONNECT: @shift_bytes 0 0 0 0 shift_bytes 0 0 0 0
-- Retrieval info: USED_PORT: status_out 0 0 8 0 OUTPUT NODEFVAL "status_out[7..0]"
-- Retrieval info: CONNECT: status_out 0 0 8 0 @status_out 0 0 8 0
-- Retrieval info: USED_PORT: write 0 0 0 0 INPUT NODEFVAL "write"
-- Retrieval info: CONNECT: @write 0 0 0 0 write 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.cmp TRUE TRUE
