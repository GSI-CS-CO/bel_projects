library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.wishbone_pkg.all;

package pwm_pkg is

    constant c_pwm_sdb : t_sdb_device := (

        abi_class     => x"0000", -- undocumented device
        abi_ver_major => x"00",
        abi_ver_minor => x"01",
        wbd_endian    => c_sdb_endian_big,
        wbd_width     => x"7", -- 8/16/32-bit port granularity
        sdb_component => (
            addr_first    => x"0000000000000000",
            addr_last     => x"0000000000000fff",
            product       => (
                vendor_id     => x"0000000000000651",
                device_id     => x"434E5453",
                version       => x"00000001",
                date          => x"20250125",
                name          => "GSI:PWM-MODULE     "
            )
        )
    );

    component pwm is

        generic (
            g_simulation                : in boolean := false;

            g_pwm_channel_num           : natural range 1 to 32 := 8;
            g_pwm_regs_size             : natural range 1 to 32 := 16;

            g_pwm_interface_mode        : t_wishbone_interface_mode := PIPELINED;
            g_pwm_address_granularity   : t_wishbone_address_granularity := BYTE
        );
        port(

            clk_sys_i       : in std_logic;
            rst_sys_n_i     : in std_logic;


            t_wb_o          : out t_wishbone_slave_out;
            t_wb_i          : in  t_wishbone_slave_in;

            pwm_latch_i     : in std_logic;
            pwm_o           : out std_logic_vector((g_pwm_channel_num-1) downto 0)
        );

    end component;

end package;