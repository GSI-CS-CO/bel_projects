LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
use work.scu_diob_pkg.all;

entity Beam_Loss_check is
    generic (
    
    WIDTH        : integer := 20     -- Counter width
       
);
port (
    clk_sys           : in std_logic;      -- Clock
    rstn_sys          : in std_logic;      -- Reset

   -- IN BLM 
    BLM_data_in       : in std_logic_vector(53 downto 0);
    BLM_gate_in       : in std_logic_vector(11 downto 0);
    BLM_tst_ck_sig    : in std_logic_vector (9 downto 0);
    --IN registers
    pos_threshold           : in t_BLM_th_Array; --t_BLM_th_Array is array (0 to 255) of std_logic_vector(31 downto 0);
    neg_threshold           : in t_BLM_th_Array ;
    BLM_wdog_hold_time_Reg  : in std_logic_vector(15 downto 0);
    BLM_gate_hold_time_Reg  : in  t_BLM_gate_hold_Time_Array;
    BLM_ctrl_Reg            : in std_logic_vector(15 downto 0); -- bit 0 = counter RESET, 
                                                                -- bit 1: when 0 the outputs of board in slot 12 are the direct outptuts of the output OR, 
                                                                --         when 1, the outputs in slot 12 are the values of AW_Output_Reg(6),   
                                                                -- bit 13..2 Direct Gate-usage, one bit for each gate signal input (BLM_gate_in), 
                                                                -- bit 14 reset from gate
                                                                -- bit 15 free

    BLM_gate_seq_ck_sel_Reg : in std_logic_vector(15 downto 0);
    BLM_gate_seq_in_ena_Reg : in std_logic_vector(15 downto 0); --"00"& ena for gate board1 &"00" & ena for gate board2 
    BLM_in_sel_Reg          : in t_BLM_reg_Array; --256 x (4 bit for gate ena & 6 bit for up signal ena & 6 for down signal ena)
    BLM_out_sel_reg : in t_BLM_out_sel_reg_Array;  --217 x 16 bits = "0000" and 6 x (54 watchdog errors+ 12 gate errors + 512 counter outputs )     

    -- OUT register
    BLM_status_Reg    : out t_IO_Reg_0_to_36_Array;
      -- OUT BLM
      BLM_Out           : out std_logic_vector(5 downto 0) 
);

end Beam_Loss_check;

architecture rtl of Beam_Loss_check is
  
  signal BLM_test_signal   : std_logic_vector(9 downto 0);  --Test signals + ground  --to reference  Test_In_Mtx
 
  signal gate_clock : std_logic_vector (11 downto 0);  
  signal g_clock: std_logic_vector(11 downto 0); 
  signal VALUE_IN:  std_logic_vector(63 downto 0);
 
  signal out_wd: std_logic_vector(53 downto 0);

  signal INT_out: std_logic_vector(53 downto 0);
  signal gate_error: std_logic_vector(11 downto 0);
  signal Gate_In_Mtx: std_logic_vector (11 downto 0):= (OTHERS => '0');  -- gate outputs from the gate timing sequence control
  signal UP_OVERFLOW: std_logic_vector(255 downto 0);     
  signal DOWN_OVERFLOW: std_logic_vector(255 downto 0);  
  signal gate_sel: integer range 0 to 255;
  signal cnt_enable: std_logic_vector(255 downto 0);
  signal BLM_Output_mtx: t_BLM_out_Array;
  signal gate_output: std_logic_vector (11 downto 0);


  component BLM_watchdog is
  
    port(
        clk_i : in std_logic;     -- chip-internal pulsed clk signal
        rstn_i : in std_logic;   -- reset signal
        hold: in std_logic_vector(15 downto 0);
        in_watchdog : in std_logic;     -- input signal
        ena_i : in std_logic;     -- enable '1' for input connected to the counter
        INTL_out: out std_logic   -- interlock output for signal that doesn't change for a given time 
    
    );
end component BLM_watchdog;

component BLM_gate_timing_seq is

    generic (
 

      n       : integer range 0 TO 12 := 12
    );
    port(
      clk_i : in std_logic_vector(n-1 downto 0);
      rstn_i : in std_logic;        -- reset signal
      gate_in : in std_logic_vector(n-1 downto 0);        -- input signal
      gate_seq_ena : in std_logic_vector(11 downto 0);     -- enable '1' for input connected to the counter
      hold_time : in  t_BLM_gate_hold_Time_Array;
      timeout_error : out std_logic_vector(n-1 downto 0); -- gate doesn't start within the given timeout
      gate_out: out std_logic_vector(n-1 downto 0)        -- out gate signal
    );
    end component BLM_gate_timing_seq;

  component  BLM_ena_in_mux is
      port (
          CLK               : in std_logic;      -- Clock
          nRST              : in std_logic;      -- Reset
          mux_sel           : in t_BLM_reg_Array;
          in_mux            : in std_logic_vector(11 downto 0);
          cnt_enable        : out std_logic_vector(255 downto 0)
      );
  end component BLM_ena_in_mux;


 component BLM_counter_pool_el is

    generic (      
        WIDTH        : integer := 20      -- Counter width
            
    );
    port (
        CLK               : in std_logic;      -- Clock
        nRST              : in std_logic;      -- Reset
        gate_reset_ena    : in std_logic;
        RESET      : in std_logic;      -- global counter reset
        ENABLE            : in std_logic;      -- Enable count operation (gate signals)
        pos_threshold     : in std_logic_vector(31 downto 0);
        neg_threshold     : in std_logic_vector(31 downto 0);
        in_counter        : in std_logic_vector(63 downto 0);
        BLM_cnt_Reg     : in std_logic_vector(15 downto 0);  -- bit 5-0 = up_in_counter select, bit 11-6 = down_in_counter select, 15..13 in_ena
        UP_OVERFLOW       : out std_logic;     -- UP_Counter overflow for the input signals
        DOWN_OVERFLOW     : out std_logic    -- DOWN_Counter overflow for the input signals

    );
  end component BLM_counter_pool_el;
  

  component  BLM_out_el is
    
      port (
        CLK              : in std_logic;      -- Clock
        nRST             : in std_logic;      -- Reset
        BLM_out_sel_reg : in t_BLM_out_sel_reg_Array;  --217 x 16 bits = "0000" and 6 x (512 counter outputs + 12 gate errors + 54 watchdog errors)                                                
      
        UP_OVERFLOW      : in std_logic_vector(255 downto 0);
        DOWN_OVERFLOW    : in std_logic_vector(255 downto 0);
      
        wd_out           : in std_logic_vector(53 downto 0); 
        gate_in          : in std_logic_vector(11 downto 0); -- to be sent to the status registers
        gate_out        : in std_logic_vector (11 downto 0); 
           
        BLM_Output      : out std_logic_vector(5 downto 0);
        BLM_status_Reg : out t_IO_Reg_0_to_36_Array
        );
     
    end component BLM_out_el;

   
---######################################################################################

begin

VALUE_IN <= BLM_test_signal & BLM_data_in;


  gate_timing_clock_sel_proc: process( BLM_gate_seq_ck_sel_Reg)
    begin
    
     for i in 0 to 11 loop
       
      

        case BLM_gate_seq_ck_sel_Reg(2 downto 0)is

          when "000" 
           =>  gate_clock(i) <= BLM_tst_ck_sig(9);  --100 MHz
          when "001" 
           =>  gate_clock(i)<= BLM_tst_ck_sig(8);   --10 MHz
          when "010" 
          =>  gate_clock(i) <= BLM_tst_ck_sig(7);   --1 MHz
          when "011" 
           =>  gate_clock (i)<= BLM_tst_ck_sig(6);   --100 kHz  
          when "100" 
           =>  gate_clock(i) <= BLM_tst_ck_sig(5);   --10 kHz
          when "101" 
           =>  gate_clock (i)<= BLM_tst_ck_sig(4);  --1 kHz
          when others 
           =>  gate_clock (i) <= NULL;
        end case;
      
 
        end loop;
    end process;

g_clock <= gate_clock;

BLM_test_signal <=  BLM_tst_ck_sig(9) & -- 100 MHz
                    BLM_tst_ck_sig(3)  & -- 99 MHz
                    BLM_tst_ck_sig(8)  & -- 10 MHz
                    BLM_tst_ck_sig(2)  & -- 9.9 MHz
                    BLM_tst_ck_sig(7)  & -- 1 MHz
                    BLM_tst_ck_sig(1)  & -- 0.99 MHz
                    BLM_tst_ck_sig(6)  & -- 100 kHz
                    BLM_tst_ck_sig(0)  & -- 99 kHz
                    BLM_tst_ck_sig(5)  & -- 10 kHz
                    '0';                 -- GND

-- for direct Gate operations: if the corresponding BLM_ctrl_Reg (bit +2)='0' then BLM_gate_in signals 
-- are used as input signal to the multiplexer  (BLM_ena_in_mux) which gives the counter enables.

direct_gate_operation: process(BLM_ctrl_Reg, BLM_gate_in, gate_output)

begin
  for i in 0 to 11 loop
    
    if BLM_ctrl_Reg(i+2) = '0' then   --when '0', gate signals are directly sent to the 12 to 256 multiplexer for the counter enables assignments
      gate_In_Mtx(i)<= BLM_gate_in(i);
    else 
      gate_IN_Mtx(i) <= gate_output(i);
    end if;
  end loop;

end process direct_gate_operation;

  gate_board: BLM_gate_timing_seq

    generic map (
      n        => 12
    )
    port map(
      clk_i => g_clock,         --
      rstn_i => rstn_sys,         -- reset signal
      gate_in => BLM_gate_in,       -- gate input signals
      gate_seq_ena => BLM_gate_seq_in_ena_Reg(13 downto 8) & BLM_gate_seq_in_ena_Reg(5 downto 0), --"00"& ena for gate board1 &"00" & ena for gate board2
      hold_time => BLM_gate_hold_time_Reg,
      timeout_error => gate_error, -- gate error
      gate_out => gate_output --gate_In_Mtx       -- out gate signal
    );
   

       wd_elem_gen: for i in 0 to 53 generate

        input_Watchdog: BLM_watchdog
         
          port map(
            clk_i => clk_sys,  
            rstn_i => rstn_sys,   -- reset signal
            hold => BLM_wdog_hold_time_Reg,
            in_watchdog => BLM_data_in(i),
            ena_i =>    '1',  -- enable for input connected to the counter
            INTL_out =>   out_wd(i));
      end generate wd_elem_gen;




---- counter ena mux ------------------------------------------------------------------------------
BLM_counter_ena_block:  BLM_ena_in_mux 
  port  map(
    CLK            => clk_sys,  
    nRST           => rstn_sys,
    mux_sel        => BLM_in_sel_Reg,
    in_mux         => gate_In_Mtx,
    cnt_enable     => cnt_enable
  );


  ---- counter pool ------------------------------------------------------------------------------

BLM_counter_pool: for i in 0 to 255 generate

BLM_counter_pool_elem: BLM_counter_pool_el
generic map (      
      WIDTH  => 20)
port map (
  CLK            => clk_sys,  
  nRST           => rstn_sys,
  gate_reset_ena => BLM_ctrl_reg(14) and cnt_enable(i),
  RESET          => BLM_ctrl_Reg(0),
  ENABLE         => cnt_enable(i),
  pos_threshold  => pos_threshold(i),
  neg_threshold  => neg_threshold(i),
  in_counter     => VALUE_IN,
  BLM_cnt_Reg    => BLM_in_sel_Reg(i),
  UP_OVERFLOW    => UP_OVERFLOW(i),
  DOWN_OVERFLOW  => DOWN_OVERFLOW(i)
  );
      end generate BLM_counter_pool;
-----------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------
-- out section


    
BLM_out_section: BLM_out_el 
     
  port map(
    CLK          => clk_sys,
    nRST           => rstn_sys,   -- Reset
    -- +++
    BLM_out_sel_reg => BLM_out_sel_reg, 
    --
    UP_OVERFLOW     => UP_OVERFLOW,
    DOWN_OVERFLOW   => DOWN_OVERFLOW,
    wd_out           => out_wd,
    gate_in         => BLM_gate_in,
    gate_out        => gate_error,
    BLM_Output      => BLM_out,
  
    BLM_status_Reg  => BLM_status_Reg 
    );

  end architecture;


