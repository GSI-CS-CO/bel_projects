altiobuf_oua_inst : altiobuf_oua PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig,
		dataout_b	 => dataout_b_sig
	);
