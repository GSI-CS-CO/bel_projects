-- megafunction wizard: %ALTREMOTE_UPDATE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altremote_update 

-- ============================================================
-- File Name: arria5_reset.vhd
-- Megafunction Name(s):
-- 			altremote_update
--
-- Simulation Library Files(s):
-- 			arriav;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altremote_update CBX_AUTO_BLACKBOX="ALL" check_app_pof="false" config_device_addr_width=32 DEVICE_FAMILY="Arria V" in_data_width=32 operation_mode="remote" out_data_width=32 busy clock data_out param read_param reconfig reset reset_timer
--VERSION_BEGIN 13.1 cbx_altremote_update 2013:10:17:04:07:49:SJ cbx_cycloneii 2013:10:17:04:07:49:SJ cbx_lpm_add_sub 2013:10:17:04:07:49:SJ cbx_lpm_compare 2013:10:17:04:07:49:SJ cbx_lpm_counter 2013:10:17:04:07:49:SJ cbx_lpm_decode 2013:10:17:04:07:49:SJ cbx_lpm_shiftreg 2013:10:17:04:07:49:SJ cbx_mgl 2013:10:17:04:34:36:SJ cbx_stratix 2013:10:17:04:07:49:SJ cbx_stratixii 2013:10:17:04:07:49:SJ  VERSION_END

 LIBRARY arriav;
 USE arriav.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = arriav_rublock 1 lpm_counter 2 reg 51 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  arria5_reset_rmtupdt_t3m IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 clock	:	IN  STD_LOGIC;
		 data_out	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 param	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 read_param	:	IN  STD_LOGIC := '0';
		 reconfig	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC;
		 reset_timer	:	IN  STD_LOGIC := '0'
	 ); 
 END arria5_reset_rmtupdt_t3m;

 ARCHITECTURE RTL OF arria5_reset_rmtupdt_t3m IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "suppress_da_rule_internal=c104;suppress_da_rule_internal=C101;suppress_da_rule_internal=C103";

	 SIGNAL	 check_busy_dffe	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe4a	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := "00000000000000000000000000000000"
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe4a_ena	:	STD_LOGIC_VECTOR(31 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe6a	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe6a_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 idle_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 idle_write_wait	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_address_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_address_state_ena	:	STD_LOGIC;
	 SIGNAL	 read_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_init_counter_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_post_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_pre_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_init_counter_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_load_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_post_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_pre_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_wait_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cntr2_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cntr3_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_sd1_regout	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w478w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w478w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w484w485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_idle524w525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable75w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rublock_regout_reg576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_range186w187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range474w492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range474w487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_all_done552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_param_start_match532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_param523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_select_shift_nloop575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w8w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_all_done536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_param_width_match537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_load496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_param522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_wait495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_range184w185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range474w475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range476w477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range479w480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_idle524w525w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address219w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address269w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address274w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address279w280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address284w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address289w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address294w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address299w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address304w305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address309w310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address314w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address224w225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address319w320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address324w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address329w330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address334w335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address229w230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address234w235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address239w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address244w245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address249w250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address254w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address259w260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address264w265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable72w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  bit_counter_all_done :	STD_LOGIC;
	 SIGNAL  bit_counter_clear :	STD_LOGIC;
	 SIGNAL  bit_counter_enable :	STD_LOGIC;
	 SIGNAL  bit_counter_param_start :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  bit_counter_param_start_match :	STD_LOGIC;
	 SIGNAL  data_in	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  idle :	STD_LOGIC;
	 SIGNAL  param_decoder_param_latch :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  param_decoder_select :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  power_up :	STD_LOGIC;
	 SIGNAL  read_address :	STD_LOGIC;
	 SIGNAL  read_data :	STD_LOGIC;
	 SIGNAL  read_init :	STD_LOGIC;
	 SIGNAL  read_init_counter :	STD_LOGIC;
	 SIGNAL  read_post :	STD_LOGIC;
	 SIGNAL  read_pre_data :	STD_LOGIC;
	 SIGNAL  rublock_captnupdt :	STD_LOGIC;
	 SIGNAL  rublock_clock :	STD_LOGIC;
	 SIGNAL  rublock_reconfig :	STD_LOGIC;
	 SIGNAL  rublock_reconfig_st :	STD_LOGIC;
	 SIGNAL  rublock_regin :	STD_LOGIC;
	 SIGNAL  rublock_regout :	STD_LOGIC;
	 SIGNAL  rublock_regout_reg :	STD_LOGIC;
	 SIGNAL  rublock_shiftnld :	STD_LOGIC;
	 SIGNAL  select_shift_nloop :	STD_LOGIC;
	 SIGNAL  shift_reg_clear :	STD_LOGIC;
	 SIGNAL  shift_reg_load_enable :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_in :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_out :	STD_LOGIC;
	 SIGNAL  shift_reg_shift_enable :	STD_LOGIC;
	 SIGNAL  start_bit_decoder_out :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  start_bit_decoder_param_select :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w22w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  w53w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  w8w :	STD_LOGIC;
	 SIGNAL  width_counter_all_done :	STD_LOGIC;
	 SIGNAL  width_counter_clear :	STD_LOGIC;
	 SIGNAL  width_counter_enable :	STD_LOGIC;
	 SIGNAL  width_counter_param_width :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  width_counter_param_width_match :	STD_LOGIC;
	 SIGNAL  width_decoder_out :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  width_decoder_param_select :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  write_data :	STD_LOGIC;
	 SIGNAL  write_init :	STD_LOGIC;
	 SIGNAL  write_init_counter :	STD_LOGIC;
	 SIGNAL  write_load :	STD_LOGIC;
	 SIGNAL  write_param	:	STD_LOGIC;
	 SIGNAL  write_post_data :	STD_LOGIC;
	 SIGNAL  write_pre_data :	STD_LOGIC;
	 SIGNAL  write_wait :	STD_LOGIC;
	 SIGNAL  wire_w_data_in_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  arriav_rublock
	 PORT
	 ( 
		captnupdt	:	IN STD_LOGIC;
		clk	:	IN STD_LOGIC;
		rconfig	:	IN STD_LOGIC;
		regin	:	IN STD_LOGIC;
		regout	:	OUT STD_LOGIC;
		rsttimer	:	IN STD_LOGIC;
		shiftnld	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w478w481w(0) <= wire_w478w(0) AND wire_w_lg_w_param_decoder_param_latch_range479w480w(0);
	wire_w_lg_w478w490w(0) <= wire_w478w(0) AND wire_w_param_decoder_param_latch_range479w(0);
	wire_w_lg_w484w485w(0) <= wire_w484w(0) AND wire_w_lg_w_param_decoder_param_latch_range479w480w(0);
	wire_w_lg_w_lg_idle524w525w(0) <= wire_w_lg_idle524w(0) AND wire_w_lg_write_param522w(0);
	wire_w493w(0) <= wire_w_lg_w_param_decoder_param_latch_range474w492w(0) AND wire_w_param_decoder_param_latch_range479w(0);
	wire_w488w(0) <= wire_w_lg_w_param_decoder_param_latch_range474w487w(0) AND wire_w_lg_w_param_decoder_param_latch_range479w480w(0);
	wire_w_lg_w_lg_read_address192w193w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range191w(0);
	wire_w_lg_w_lg_read_address192w228w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range227w(0);
	wire_w_lg_w_lg_read_address192w233w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range232w(0);
	wire_w_lg_w_lg_read_address192w238w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range237w(0);
	wire_w_lg_w_lg_read_address192w243w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range242w(0);
	wire_w_lg_w_lg_read_address192w248w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range247w(0);
	wire_w_lg_w_lg_read_address192w253w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range252w(0);
	wire_w_lg_w_lg_read_address192w258w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range257w(0);
	wire_w_lg_w_lg_read_address192w263w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range262w(0);
	wire_w_lg_w_lg_read_address192w268w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range267w(0);
	wire_w_lg_w_lg_read_address192w273w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range272w(0);
	wire_w_lg_w_lg_read_address192w197w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range196w(0);
	wire_w_lg_w_lg_read_address192w278w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range277w(0);
	wire_w_lg_w_lg_read_address192w283w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range282w(0);
	wire_w_lg_w_lg_read_address192w288w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range287w(0);
	wire_w_lg_w_lg_read_address192w293w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range292w(0);
	wire_w_lg_w_lg_read_address192w298w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range297w(0);
	wire_w_lg_w_lg_read_address192w303w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range302w(0);
	wire_w_lg_w_lg_read_address192w308w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range307w(0);
	wire_w_lg_w_lg_read_address192w313w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range312w(0);
	wire_w_lg_w_lg_read_address192w318w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range317w(0);
	wire_w_lg_w_lg_read_address192w323w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range322w(0);
	wire_w_lg_w_lg_read_address192w200w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range199w(0);
	wire_w_lg_w_lg_read_address192w328w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range327w(0);
	wire_w_lg_w_lg_read_address192w333w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range332w(0);
	wire_w_lg_w_lg_read_address192w203w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range202w(0);
	wire_w_lg_w_lg_read_address192w206w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range205w(0);
	wire_w_lg_w_lg_read_address192w209w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range208w(0);
	wire_w_lg_w_lg_read_address192w212w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range211w(0);
	wire_w_lg_w_lg_read_address192w215w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range214w(0);
	wire_w_lg_w_lg_read_address192w218w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range217w(0);
	wire_w_lg_w_lg_read_address192w223w(0) <= wire_w_lg_read_address192w(0) AND wire_dffe4a_w_q_range222w(0);
	wire_w_lg_w_lg_shift_reg_load_enable75w77w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(1);
	wire_w_lg_w_lg_shift_reg_load_enable75w113w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(10);
	wire_w_lg_w_lg_shift_reg_load_enable75w117w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(11);
	wire_w_lg_w_lg_shift_reg_load_enable75w121w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(12);
	wire_w_lg_w_lg_shift_reg_load_enable75w125w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(13);
	wire_w_lg_w_lg_shift_reg_load_enable75w129w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(14);
	wire_w_lg_w_lg_shift_reg_load_enable75w133w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(15);
	wire_w_lg_w_lg_shift_reg_load_enable75w137w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(16);
	wire_w_lg_w_lg_shift_reg_load_enable75w141w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(17);
	wire_w_lg_w_lg_shift_reg_load_enable75w145w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(18);
	wire_w_lg_w_lg_shift_reg_load_enable75w149w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(19);
	wire_w_lg_w_lg_shift_reg_load_enable75w81w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(2);
	wire_w_lg_w_lg_shift_reg_load_enable75w153w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(20);
	wire_w_lg_w_lg_shift_reg_load_enable75w157w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(21);
	wire_w_lg_w_lg_shift_reg_load_enable75w161w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(22);
	wire_w_lg_w_lg_shift_reg_load_enable75w165w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(23);
	wire_w_lg_w_lg_shift_reg_load_enable75w169w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(24);
	wire_w_lg_w_lg_shift_reg_load_enable75w85w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(3);
	wire_w_lg_w_lg_shift_reg_load_enable75w89w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(4);
	wire_w_lg_w_lg_shift_reg_load_enable75w93w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(5);
	wire_w_lg_w_lg_shift_reg_load_enable75w97w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(6);
	wire_w_lg_w_lg_shift_reg_load_enable75w101w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(7);
	wire_w_lg_w_lg_shift_reg_load_enable75w105w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(8);
	wire_w_lg_w_lg_shift_reg_load_enable75w109w(0) <= wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(9);
	wire_w478w(0) <= wire_w_lg_w_param_decoder_param_latch_range474w475w(0) AND wire_w_lg_w_param_decoder_param_latch_range476w477w(0);
	wire_w484w(0) <= wire_w_lg_w_param_decoder_param_latch_range474w475w(0) AND wire_w_param_decoder_param_latch_range476w(0);
	wire_w_lg_idle524w(0) <= idle AND wire_w_lg_read_param523w(0);
	wire_w_lg_read_address219w(0) <= read_address AND wire_dffe4a_w_q_range191w(0);
	wire_w_lg_read_address269w(0) <= read_address AND wire_dffe4a_w_q_range227w(0);
	wire_w_lg_read_address274w(0) <= read_address AND wire_dffe4a_w_q_range232w(0);
	wire_w_lg_read_address279w(0) <= read_address AND wire_dffe4a_w_q_range237w(0);
	wire_w_lg_read_address284w(0) <= read_address AND wire_dffe4a_w_q_range242w(0);
	wire_w_lg_read_address289w(0) <= read_address AND wire_dffe4a_w_q_range247w(0);
	wire_w_lg_read_address294w(0) <= read_address AND wire_dffe4a_w_q_range252w(0);
	wire_w_lg_read_address299w(0) <= read_address AND wire_dffe4a_w_q_range257w(0);
	wire_w_lg_read_address304w(0) <= read_address AND wire_dffe4a_w_q_range262w(0);
	wire_w_lg_read_address309w(0) <= read_address AND wire_dffe4a_w_q_range267w(0);
	wire_w_lg_read_address314w(0) <= read_address AND wire_dffe4a_w_q_range272w(0);
	wire_w_lg_read_address224w(0) <= read_address AND wire_dffe4a_w_q_range196w(0);
	wire_w_lg_read_address319w(0) <= read_address AND wire_dffe4a_w_q_range277w(0);
	wire_w_lg_read_address324w(0) <= read_address AND wire_dffe4a_w_q_range282w(0);
	wire_w_lg_read_address329w(0) <= read_address AND wire_dffe4a_w_q_range287w(0);
	wire_w_lg_read_address334w(0) <= read_address AND wire_dffe4a_w_q_range292w(0);
	wire_w_lg_read_address229w(0) <= read_address AND wire_dffe4a_w_q_range199w(0);
	wire_w_lg_read_address234w(0) <= read_address AND wire_dffe4a_w_q_range202w(0);
	wire_w_lg_read_address239w(0) <= read_address AND wire_dffe4a_w_q_range205w(0);
	wire_w_lg_read_address244w(0) <= read_address AND wire_dffe4a_w_q_range208w(0);
	wire_w_lg_read_address249w(0) <= read_address AND wire_dffe4a_w_q_range211w(0);
	wire_w_lg_read_address254w(0) <= read_address AND wire_dffe4a_w_q_range214w(0);
	wire_w_lg_read_address259w(0) <= read_address AND wire_dffe4a_w_q_range217w(0);
	wire_w_lg_read_address264w(0) <= read_address AND wire_dffe4a_w_q_range222w(0);
	wire_w_lg_read_data538w(0) <= read_data AND wire_w_lg_width_counter_param_width_match537w(0);
	wire_w_lg_read_init_counter534w(0) <= read_init_counter AND wire_w_lg_bit_counter_param_start_match532w(0);
	wire_w_lg_read_post544w(0) <= read_post AND wire_w_lg_width_counter_all_done536w(0);
	wire_w_lg_read_pre_data533w(0) <= read_pre_data AND wire_w_lg_bit_counter_param_start_match532w(0);
	wire_w_lg_rublock_regout_reg576w(0) <= rublock_regout_reg AND wire_w_lg_select_shift_nloop575w(0);
	wire_w_lg_shift_reg_load_enable87w(0) <= shift_reg_load_enable AND wire_w_data_in_range86w(0);
	wire_w_lg_shift_reg_load_enable91w(0) <= shift_reg_load_enable AND wire_w_data_in_range90w(0);
	wire_w_lg_shift_reg_load_enable95w(0) <= shift_reg_load_enable AND wire_w_data_in_range94w(0);
	wire_w_lg_shift_reg_load_enable99w(0) <= shift_reg_load_enable AND wire_w_data_in_range98w(0);
	wire_w_lg_shift_reg_load_enable103w(0) <= shift_reg_load_enable AND wire_w_data_in_range102w(0);
	wire_w_lg_shift_reg_load_enable107w(0) <= shift_reg_load_enable AND wire_w_data_in_range106w(0);
	wire_w_lg_shift_reg_load_enable111w(0) <= shift_reg_load_enable AND wire_w_data_in_range110w(0);
	wire_w_lg_shift_reg_load_enable115w(0) <= shift_reg_load_enable AND wire_w_data_in_range114w(0);
	wire_w_lg_shift_reg_load_enable119w(0) <= shift_reg_load_enable AND wire_w_data_in_range118w(0);
	wire_w_lg_shift_reg_load_enable123w(0) <= shift_reg_load_enable AND wire_w_data_in_range122w(0);
	wire_w_lg_shift_reg_load_enable127w(0) <= shift_reg_load_enable AND wire_w_data_in_range126w(0);
	wire_w_lg_shift_reg_load_enable131w(0) <= shift_reg_load_enable AND wire_w_data_in_range130w(0);
	wire_w_lg_shift_reg_load_enable135w(0) <= shift_reg_load_enable AND wire_w_data_in_range134w(0);
	wire_w_lg_shift_reg_load_enable139w(0) <= shift_reg_load_enable AND wire_w_data_in_range138w(0);
	wire_w_lg_shift_reg_load_enable143w(0) <= shift_reg_load_enable AND wire_w_data_in_range142w(0);
	wire_w_lg_shift_reg_load_enable147w(0) <= shift_reg_load_enable AND wire_w_data_in_range146w(0);
	wire_w_lg_shift_reg_load_enable151w(0) <= shift_reg_load_enable AND wire_w_data_in_range150w(0);
	wire_w_lg_shift_reg_load_enable155w(0) <= shift_reg_load_enable AND wire_w_data_in_range154w(0);
	wire_w_lg_shift_reg_load_enable159w(0) <= shift_reg_load_enable AND wire_w_data_in_range158w(0);
	wire_w_lg_shift_reg_load_enable163w(0) <= shift_reg_load_enable AND wire_w_data_in_range162w(0);
	wire_w_lg_shift_reg_load_enable167w(0) <= shift_reg_load_enable AND wire_w_data_in_range166w(0);
	wire_w_lg_shift_reg_load_enable171w(0) <= shift_reg_load_enable AND wire_w_data_in_range170w(0);
	wire_w_lg_shift_reg_load_enable79w(0) <= shift_reg_load_enable AND wire_w_data_in_range78w(0);
	wire_w_lg_shift_reg_load_enable83w(0) <= shift_reg_load_enable AND wire_w_data_in_range82w(0);
	wire_w_lg_write_data553w(0) <= write_data AND wire_w_lg_width_counter_param_width_match537w(0);
	wire_w_lg_write_init_counter550w(0) <= write_init_counter AND wire_w_lg_bit_counter_param_start_match532w(0);
	wire_w_lg_write_post_data559w(0) <= write_post_data AND wire_w_lg_bit_counter_all_done552w(0);
	wire_w_lg_write_pre_data549w(0) <= write_pre_data AND wire_w_lg_bit_counter_param_start_match532w(0);
	wire_w_lg_w_param_range186w187w(0) <= wire_w_param_range186w(0) AND wire_w_lg_w_param_range184w185w(0);
	wire_w_lg_w_param_decoder_param_latch_range474w492w(0) <= wire_w_param_decoder_param_latch_range474w(0) AND wire_w_lg_w_param_decoder_param_latch_range476w477w(0);
	wire_w_lg_w_param_decoder_param_latch_range474w487w(0) <= wire_w_param_decoder_param_latch_range474w(0) AND wire_w_param_decoder_param_latch_range476w(0);
	wire_w_lg_bit_counter_all_done552w(0) <= NOT bit_counter_all_done;
	wire_w_lg_bit_counter_param_start_match532w(0) <= NOT bit_counter_param_start_match;
	wire_w_lg_idle507w(0) <= NOT idle;
	wire_w_lg_read_address192w(0) <= NOT read_address;
	wire_w_lg_read_data503w(0) <= NOT read_data;
	wire_w_lg_read_init506w(0) <= NOT read_init;
	wire_w_lg_read_init_counter505w(0) <= NOT read_init_counter;
	wire_w_lg_read_param523w(0) <= NOT read_param;
	wire_w_lg_read_post502w(0) <= NOT read_post;
	wire_w_lg_read_pre_data504w(0) <= NOT read_pre_data;
	wire_w_lg_select_shift_nloop575w(0) <= NOT select_shift_nloop;
	wire_w_lg_shift_reg_load_enable75w(0) <= NOT shift_reg_load_enable;
	wire_w_lg_w8w181w(0) <= NOT w8w;
	wire_w_lg_width_counter_all_done536w(0) <= NOT width_counter_all_done;
	wire_w_lg_width_counter_param_width_match537w(0) <= NOT width_counter_param_width_match;
	wire_w_lg_write_data498w(0) <= NOT write_data;
	wire_w_lg_write_init501w(0) <= NOT write_init;
	wire_w_lg_write_init_counter500w(0) <= NOT write_init_counter;
	wire_w_lg_write_load496w(0) <= NOT write_load;
	wire_w_lg_write_param522w(0) <= NOT write_param;
	wire_w_lg_write_post_data497w(0) <= NOT write_post_data;
	wire_w_lg_write_pre_data499w(0) <= NOT write_pre_data;
	wire_w_lg_write_wait495w(0) <= NOT write_wait;
	wire_w_lg_w_param_range184w185w(0) <= NOT wire_w_param_range184w(0);
	wire_w_lg_w_param_decoder_param_latch_range474w475w(0) <= NOT wire_w_param_decoder_param_latch_range474w(0);
	wire_w_lg_w_param_decoder_param_latch_range476w477w(0) <= NOT wire_w_param_decoder_param_latch_range476w(0);
	wire_w_lg_w_param_decoder_param_latch_range479w480w(0) <= NOT wire_w_param_decoder_param_latch_range479w(0);
	wire_w_lg_w_lg_w_lg_idle524w525w526w(0) <= wire_w_lg_w_lg_idle524w525w(0) OR write_wait;
	wire_w_lg_w_lg_read_address219w220w(0) <= wire_w_lg_read_address219w(0) OR wire_w_lg_w_lg_read_address192w218w(0);
	wire_w_lg_w_lg_read_address269w270w(0) <= wire_w_lg_read_address269w(0) OR wire_w_lg_w_lg_read_address192w268w(0);
	wire_w_lg_w_lg_read_address274w275w(0) <= wire_w_lg_read_address274w(0) OR wire_w_lg_w_lg_read_address192w273w(0);
	wire_w_lg_w_lg_read_address279w280w(0) <= wire_w_lg_read_address279w(0) OR wire_w_lg_w_lg_read_address192w278w(0);
	wire_w_lg_w_lg_read_address284w285w(0) <= wire_w_lg_read_address284w(0) OR wire_w_lg_w_lg_read_address192w283w(0);
	wire_w_lg_w_lg_read_address289w290w(0) <= wire_w_lg_read_address289w(0) OR wire_w_lg_w_lg_read_address192w288w(0);
	wire_w_lg_w_lg_read_address294w295w(0) <= wire_w_lg_read_address294w(0) OR wire_w_lg_w_lg_read_address192w293w(0);
	wire_w_lg_w_lg_read_address299w300w(0) <= wire_w_lg_read_address299w(0) OR wire_w_lg_w_lg_read_address192w298w(0);
	wire_w_lg_w_lg_read_address304w305w(0) <= wire_w_lg_read_address304w(0) OR wire_w_lg_w_lg_read_address192w303w(0);
	wire_w_lg_w_lg_read_address309w310w(0) <= wire_w_lg_read_address309w(0) OR wire_w_lg_w_lg_read_address192w308w(0);
	wire_w_lg_w_lg_read_address314w315w(0) <= wire_w_lg_read_address314w(0) OR wire_w_lg_w_lg_read_address192w313w(0);
	wire_w_lg_w_lg_read_address224w225w(0) <= wire_w_lg_read_address224w(0) OR wire_w_lg_w_lg_read_address192w223w(0);
	wire_w_lg_w_lg_read_address319w320w(0) <= wire_w_lg_read_address319w(0) OR wire_w_lg_w_lg_read_address192w318w(0);
	wire_w_lg_w_lg_read_address324w325w(0) <= wire_w_lg_read_address324w(0) OR wire_w_lg_w_lg_read_address192w323w(0);
	wire_w_lg_w_lg_read_address329w330w(0) <= wire_w_lg_read_address329w(0) OR wire_w_lg_w_lg_read_address192w328w(0);
	wire_w_lg_w_lg_read_address334w335w(0) <= wire_w_lg_read_address334w(0) OR wire_w_lg_w_lg_read_address192w333w(0);
	wire_w_lg_w_lg_read_address229w230w(0) <= wire_w_lg_read_address229w(0) OR wire_w_lg_w_lg_read_address192w228w(0);
	wire_w_lg_w_lg_read_address234w235w(0) <= wire_w_lg_read_address234w(0) OR wire_w_lg_w_lg_read_address192w233w(0);
	wire_w_lg_w_lg_read_address239w240w(0) <= wire_w_lg_read_address239w(0) OR wire_w_lg_w_lg_read_address192w238w(0);
	wire_w_lg_w_lg_read_address244w245w(0) <= wire_w_lg_read_address244w(0) OR wire_w_lg_w_lg_read_address192w243w(0);
	wire_w_lg_w_lg_read_address249w250w(0) <= wire_w_lg_read_address249w(0) OR wire_w_lg_w_lg_read_address192w248w(0);
	wire_w_lg_w_lg_read_address254w255w(0) <= wire_w_lg_read_address254w(0) OR wire_w_lg_w_lg_read_address192w253w(0);
	wire_w_lg_w_lg_read_address259w260w(0) <= wire_w_lg_read_address259w(0) OR wire_w_lg_w_lg_read_address192w258w(0);
	wire_w_lg_w_lg_read_address264w265w(0) <= wire_w_lg_read_address264w(0) OR wire_w_lg_w_lg_read_address192w263w(0);
	wire_w_lg_w_lg_shift_reg_load_enable72w73w(0) <= wire_w_lg_shift_reg_load_enable72w(0) OR shift_reg_clear;
	wire_w_lg_shift_reg_load_enable72w(0) <= shift_reg_load_enable OR shift_reg_shift_enable;
	bit_counter_all_done <= (((((wire_cntr2_q(0) AND wire_cntr2_q(1)) AND (NOT wire_cntr2_q(2))) AND wire_cntr2_q(3)) AND (NOT wire_cntr2_q(4))) AND wire_cntr2_q(5));
	bit_counter_clear <= (read_init OR write_init);
	bit_counter_enable <= (((((((((read_init OR write_init) OR read_init_counter) OR write_init_counter) OR read_pre_data) OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data);
	bit_counter_param_start <= start_bit_decoder_out;
	bit_counter_param_start_match <= ((((((NOT w22w(0)) AND (NOT w22w(1))) AND (NOT w22w(2))) AND (NOT w22w(3))) AND (NOT w22w(4))) AND (NOT w22w(5)));
	busy <= wire_w_lg_idle507w(0);
	data_in <= (OTHERS => '0');
	data_out <= ( wire_w_lg_w_lg_read_address334w335w & wire_w_lg_w_lg_read_address329w330w & wire_w_lg_w_lg_read_address324w325w & wire_w_lg_w_lg_read_address319w320w & wire_w_lg_w_lg_read_address314w315w & wire_w_lg_w_lg_read_address309w310w & wire_w_lg_w_lg_read_address304w305w & wire_w_lg_w_lg_read_address299w300w & wire_w_lg_w_lg_read_address294w295w & wire_w_lg_w_lg_read_address289w290w & wire_w_lg_w_lg_read_address284w285w & wire_w_lg_w_lg_read_address279w280w & wire_w_lg_w_lg_read_address274w275w & wire_w_lg_w_lg_read_address269w270w & wire_w_lg_w_lg_read_address264w265w & wire_w_lg_w_lg_read_address259w260w & wire_w_lg_w_lg_read_address254w255w & wire_w_lg_w_lg_read_address249w250w & wire_w_lg_w_lg_read_address244w245w & wire_w_lg_w_lg_read_address239w240w & wire_w_lg_w_lg_read_address234w235w & wire_w_lg_w_lg_read_address229w230w & wire_w_lg_w_lg_read_address224w225w & wire_w_lg_w_lg_read_address219w220w & wire_w_lg_w_lg_read_address192w215w & wire_w_lg_w_lg_read_address192w212w & wire_w_lg_w_lg_read_address192w209w & wire_w_lg_w_lg_read_address192w206w & wire_w_lg_w_lg_read_address192w203w & wire_w_lg_w_lg_read_address192w200w & wire_w_lg_w_lg_read_address192w197w & wire_w_lg_w_lg_read_address192w193w);
	idle <= idle_state;
	param_decoder_param_latch <= dffe6a;
	param_decoder_select <= ( wire_w493w & wire_w_lg_w478w490w & wire_w488w & wire_w_lg_w484w485w & wire_w_lg_w478w481w);
	power_up <= ((((((((((((wire_w_lg_idle507w(0) AND wire_w_lg_read_init506w(0)) AND wire_w_lg_read_init_counter505w(0)) AND wire_w_lg_read_pre_data504w(0)) AND wire_w_lg_read_data503w(0)) AND wire_w_lg_read_post502w(0)) AND wire_w_lg_write_init501w(0)) AND wire_w_lg_write_init_counter500w(0)) AND wire_w_lg_write_pre_data499w(0)) AND wire_w_lg_write_data498w(0)) AND wire_w_lg_write_post_data497w(0)) AND wire_w_lg_write_load496w(0)) AND wire_w_lg_write_wait495w(0));
	read_address <= read_address_state;
	read_data <= read_data_state;
	read_init <= read_init_state;
	read_init_counter <= read_init_counter_state;
	read_post <= read_post_state;
	read_pre_data <= read_pre_data_state;
	rublock_captnupdt <= wire_w_lg_write_load496w(0);
	rublock_clock <= (NOT (clock OR idle_write_wait));
	rublock_reconfig <= rublock_reconfig_st;
	rublock_reconfig_st <= (idle AND reconfig);
	rublock_regin <= (wire_w_lg_rublock_regout_reg576w(0) OR (shift_reg_serial_out AND select_shift_nloop));
	rublock_regout <= wire_sd1_regout;
	rublock_regout_reg <= dffe5;
	rublock_shiftnld <= (((((read_pre_data OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data);
	select_shift_nloop <= (wire_w_lg_read_data538w(0) OR wire_w_lg_write_data553w(0));
	shift_reg_clear <= read_init;
	shift_reg_load_enable <= (idle AND write_param);
	shift_reg_serial_in <= (rublock_regout_reg AND select_shift_nloop);
	shift_reg_serial_out <= dffe4a(0);
	shift_reg_shift_enable <= (((read_data OR write_data) OR read_post) OR write_post_data);
	start_bit_decoder_out <= ((((( "0" & "0" & "0" & "0" & "0" & "0") OR ( "0" & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1))) OR ( "0" & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & "0")) OR ( "0" & "0" & "0" & start_bit_decoder_param_select(3) & start_bit_decoder_param_select(3) & "0")) OR ( "0" & "0" & "0" & start_bit_decoder_param_select(4) & "0" & start_bit_decoder_param_select(4)));
	start_bit_decoder_param_select <= param_decoder_select;
	w22w <= (wire_cntr2_q XOR bit_counter_param_start);
	w53w <= (wire_cntr3_q XOR width_counter_param_width);
	w8w <= wire_w_lg_idle507w(0);
	width_counter_all_done <= (((((wire_cntr3_q(0) AND wire_cntr3_q(1)) AND wire_cntr3_q(2)) AND wire_cntr3_q(3)) AND wire_cntr3_q(4)) AND (NOT wire_cntr3_q(5)));
	width_counter_clear <= (read_init OR write_init);
	width_counter_enable <= ((read_data OR write_data) OR read_post);
	width_counter_param_width <= width_decoder_out;
	width_counter_param_width_match <= ((((((NOT w53w(0)) AND (NOT w53w(1))) AND (NOT w53w(2))) AND (NOT w53w(3))) AND (NOT w53w(4))) AND (NOT w53w(5)));
	width_decoder_out <= ((((( "0" & "0" & "0" & width_decoder_param_select(0) & "0" & width_decoder_param_select(0)) OR ( "0" & "0" & width_decoder_param_select(1) & width_decoder_param_select(1) & "0" & "0")) OR ( "0" & "0" & "0" & "0" & "0" & width_decoder_param_select(2))) OR ( "0" & width_decoder_param_select(3) & width_decoder_param_select(3) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & "0" & "0" & width_decoder_param_select(4)));
	width_decoder_param_select <= param_decoder_select;
	write_data <= write_data_state;
	write_init <= write_init_state;
	write_init_counter <= write_init_counter_state;
	write_load <= write_load_state;
	write_param <= '0';
	write_post_data <= write_post_data_state;
	write_pre_data <= write_pre_data_state;
	write_wait <= write_wait_state;
	wire_w_data_in_range86w(0) <= data_in(10);
	wire_w_data_in_range90w(0) <= data_in(11);
	wire_w_data_in_range94w(0) <= data_in(12);
	wire_w_data_in_range98w(0) <= data_in(13);
	wire_w_data_in_range102w(0) <= data_in(14);
	wire_w_data_in_range106w(0) <= data_in(15);
	wire_w_data_in_range110w(0) <= data_in(16);
	wire_w_data_in_range114w(0) <= data_in(17);
	wire_w_data_in_range118w(0) <= data_in(18);
	wire_w_data_in_range122w(0) <= data_in(19);
	wire_w_data_in_range126w(0) <= data_in(20);
	wire_w_data_in_range130w(0) <= data_in(21);
	wire_w_data_in_range134w(0) <= data_in(22);
	wire_w_data_in_range138w(0) <= data_in(23);
	wire_w_data_in_range142w(0) <= data_in(24);
	wire_w_data_in_range146w(0) <= data_in(25);
	wire_w_data_in_range150w(0) <= data_in(26);
	wire_w_data_in_range154w(0) <= data_in(27);
	wire_w_data_in_range158w(0) <= data_in(28);
	wire_w_data_in_range162w(0) <= data_in(29);
	wire_w_data_in_range166w(0) <= data_in(30);
	wire_w_data_in_range170w(0) <= data_in(31);
	wire_w_data_in_range78w(0) <= data_in(8);
	wire_w_data_in_range82w(0) <= data_in(9);
	wire_w_param_range184w(0) <= param(1);
	wire_w_param_range186w(0) <= param(2);
	wire_w_param_decoder_param_latch_range474w(0) <= param_decoder_param_latch(0);
	wire_w_param_decoder_param_latch_range476w(0) <= param_decoder_param_latch(1);
	wire_w_param_decoder_param_latch_range479w(0) <= param_decoder_param_latch(2);
	check_busy_dffe <= (OTHERS => '0');
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(0) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(0) <= '0';
				ELSE dffe4a(0) <= (wire_w_lg_shift_reg_load_enable79w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w77w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(1) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(1) <= '0';
				ELSE dffe4a(1) <= (wire_w_lg_shift_reg_load_enable83w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w81w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(2) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(2) <= '0';
				ELSE dffe4a(2) <= (wire_w_lg_shift_reg_load_enable87w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w85w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(3) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(3) <= '0';
				ELSE dffe4a(3) <= (wire_w_lg_shift_reg_load_enable91w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w89w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(4) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(4) <= '0';
				ELSE dffe4a(4) <= (wire_w_lg_shift_reg_load_enable95w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w93w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(5) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(5) <= '0';
				ELSE dffe4a(5) <= (wire_w_lg_shift_reg_load_enable99w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w97w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(6) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(6) <= '0';
				ELSE dffe4a(6) <= (wire_w_lg_shift_reg_load_enable103w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w101w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(7) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(7) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(7) <= '0';
				ELSE dffe4a(7) <= (wire_w_lg_shift_reg_load_enable107w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w105w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(8) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(8) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(8) <= '0';
				ELSE dffe4a(8) <= (wire_w_lg_shift_reg_load_enable111w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w109w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(9) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(9) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(9) <= '0';
				ELSE dffe4a(9) <= (wire_w_lg_shift_reg_load_enable115w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w113w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(10) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(10) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(10) <= '0';
				ELSE dffe4a(10) <= (wire_w_lg_shift_reg_load_enable119w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w117w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(11) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(11) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(11) <= '0';
				ELSE dffe4a(11) <= (wire_w_lg_shift_reg_load_enable123w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w121w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(12) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(12) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(12) <= '0';
				ELSE dffe4a(12) <= (wire_w_lg_shift_reg_load_enable127w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w125w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(13) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(13) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(13) <= '0';
				ELSE dffe4a(13) <= (wire_w_lg_shift_reg_load_enable131w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w129w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(14) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(14) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(14) <= '0';
				ELSE dffe4a(14) <= (wire_w_lg_shift_reg_load_enable135w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w133w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(15) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(15) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(15) <= '0';
				ELSE dffe4a(15) <= (wire_w_lg_shift_reg_load_enable139w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w137w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(16) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(16) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(16) <= '0';
				ELSE dffe4a(16) <= (wire_w_lg_shift_reg_load_enable143w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w141w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(17) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(17) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(17) <= '0';
				ELSE dffe4a(17) <= (wire_w_lg_shift_reg_load_enable147w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w145w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(18) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(18) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(18) <= '0';
				ELSE dffe4a(18) <= (wire_w_lg_shift_reg_load_enable151w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w149w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(19) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(19) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(19) <= '0';
				ELSE dffe4a(19) <= (wire_w_lg_shift_reg_load_enable155w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w153w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(20) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(20) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(20) <= '0';
				ELSE dffe4a(20) <= (wire_w_lg_shift_reg_load_enable159w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w157w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(21) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(21) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(21) <= '0';
				ELSE dffe4a(21) <= (wire_w_lg_shift_reg_load_enable163w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w161w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(22) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(22) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(22) <= '0';
				ELSE dffe4a(22) <= (wire_w_lg_shift_reg_load_enable167w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w165w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(23) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(23) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(23) <= '0';
				ELSE dffe4a(23) <= (wire_w_lg_shift_reg_load_enable171w(0) OR wire_w_lg_w_lg_shift_reg_load_enable75w169w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(24) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(24) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(24) <= '0';
				ELSE dffe4a(24) <= (wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(25));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(25) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(25) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(25) <= '0';
				ELSE dffe4a(25) <= (wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(26));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(26) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(26) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(26) <= '0';
				ELSE dffe4a(26) <= (wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(27));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(27) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(27) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(27) <= '0';
				ELSE dffe4a(27) <= (wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(28));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(28) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(28) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(28) <= '0';
				ELSE dffe4a(28) <= (wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(29));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(29) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(29) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(29) <= '0';
				ELSE dffe4a(29) <= (wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(30));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(30) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(30) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(30) <= '0';
				ELSE dffe4a(30) <= (wire_w_lg_shift_reg_load_enable75w(0) AND dffe4a(31));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(31) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(31) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(31) <= '0';
				ELSE dffe4a(31) <= (wire_w_lg_shift_reg_load_enable75w(0) AND shift_reg_serial_in);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	loop0 : FOR i IN 0 TO 31 GENERATE
		wire_dffe4a_ena(i) <= wire_w_lg_w_lg_shift_reg_load_enable72w73w(0);
	END GENERATE loop0;
	wire_dffe4a_w_q_range191w(0) <= dffe4a(0);
	wire_dffe4a_w_q_range227w(0) <= dffe4a(10);
	wire_dffe4a_w_q_range232w(0) <= dffe4a(11);
	wire_dffe4a_w_q_range237w(0) <= dffe4a(12);
	wire_dffe4a_w_q_range242w(0) <= dffe4a(13);
	wire_dffe4a_w_q_range247w(0) <= dffe4a(14);
	wire_dffe4a_w_q_range252w(0) <= dffe4a(15);
	wire_dffe4a_w_q_range257w(0) <= dffe4a(16);
	wire_dffe4a_w_q_range262w(0) <= dffe4a(17);
	wire_dffe4a_w_q_range267w(0) <= dffe4a(18);
	wire_dffe4a_w_q_range272w(0) <= dffe4a(19);
	wire_dffe4a_w_q_range196w(0) <= dffe4a(1);
	wire_dffe4a_w_q_range277w(0) <= dffe4a(20);
	wire_dffe4a_w_q_range282w(0) <= dffe4a(21);
	wire_dffe4a_w_q_range287w(0) <= dffe4a(22);
	wire_dffe4a_w_q_range292w(0) <= dffe4a(23);
	wire_dffe4a_w_q_range297w(0) <= dffe4a(24);
	wire_dffe4a_w_q_range302w(0) <= dffe4a(25);
	wire_dffe4a_w_q_range307w(0) <= dffe4a(26);
	wire_dffe4a_w_q_range312w(0) <= dffe4a(27);
	wire_dffe4a_w_q_range317w(0) <= dffe4a(28);
	wire_dffe4a_w_q_range322w(0) <= dffe4a(29);
	wire_dffe4a_w_q_range199w(0) <= dffe4a(2);
	wire_dffe4a_w_q_range327w(0) <= dffe4a(30);
	wire_dffe4a_w_q_range332w(0) <= dffe4a(31);
	wire_dffe4a_w_q_range202w(0) <= dffe4a(3);
	wire_dffe4a_w_q_range205w(0) <= dffe4a(4);
	wire_dffe4a_w_q_range208w(0) <= dffe4a(5);
	wire_dffe4a_w_q_range211w(0) <= dffe4a(6);
	wire_dffe4a_w_q_range214w(0) <= dffe4a(7);
	wire_dffe4a_w_q_range217w(0) <= dffe4a(8);
	wire_dffe4a_w_q_range222w(0) <= dffe4a(9);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe5 <= rublock_regout;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe6a(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe6a_ena(0) = '1') THEN dffe6a(0) <= param(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe6a(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe6a_ena(1) = '1') THEN dffe6a(1) <= param(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe6a(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe6a_ena(2) = '1') THEN dffe6a(2) <= param(2);
			END IF;
		END IF;
	END PROCESS;
	loop1 : FOR i IN 0 TO 2 GENERATE
		wire_dffe6a_ena(i) <= (idle AND (write_param OR read_param));
	END GENERATE loop1;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN idle_state <= '1';
		ELSIF (clock = '1' AND clock'event) THEN idle_state <= (((wire_w_lg_w_lg_w_lg_idle524w525w526w(0) OR (read_data AND width_counter_all_done)) OR (read_post AND width_counter_all_done)) OR power_up);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN idle_write_wait <= '0';
		ELSIF (clock = '1' AND clock'event) THEN idle_write_wait <= ((((wire_w_lg_w_lg_w_lg_idle524w525w526w(0) OR (read_data AND width_counter_all_done)) OR (read_post AND width_counter_all_done)) OR power_up) AND write_load);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_address_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_read_address_state_ena = '1') THEN read_address_state <= (((read_param OR write_param) AND (wire_w_lg_w_param_range186w187w(0) AND (NOT param(0)))) AND wire_w_lg_w8w181w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_read_address_state_ena <= (read_param OR write_param);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_data_state <= (((read_init_counter AND bit_counter_param_start_match) OR (read_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_read_data538w(0) AND wire_w_lg_width_counter_all_done536w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_init_counter_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_init_counter_state <= read_init;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_init_state <= (idle AND read_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_post_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_post_state <= (((read_data AND width_counter_param_width_match) AND wire_w_lg_width_counter_all_done536w(0)) OR wire_w_lg_read_post544w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_pre_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_pre_data_state <= (wire_w_lg_read_init_counter534w(0) OR wire_w_lg_read_pre_data533w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_data_state <= (((write_init_counter AND bit_counter_param_start_match) OR (write_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_write_data553w(0) AND wire_w_lg_bit_counter_all_done552w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_init_counter_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_init_counter_state <= write_init;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_init_state <= (idle AND write_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_load_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_load_state <= ((write_data AND bit_counter_all_done) OR (write_post_data AND bit_counter_all_done));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_post_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_post_data_state <= (((write_data AND width_counter_param_width_match) AND wire_w_lg_bit_counter_all_done552w(0)) OR wire_w_lg_write_post_data559w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_pre_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_pre_data_state <= (wire_w_lg_write_init_counter550w(0) OR wire_w_lg_write_pre_data549w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_wait_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_wait_state <= write_load;
		END IF;
	END PROCESS;
	cntr2 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		aclr => reset,
		clock => clock,
		cnt_en => bit_counter_enable,
		q => wire_cntr2_q,
		sclr => bit_counter_clear
	  );
	cntr3 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		aclr => reset,
		clock => clock,
		cnt_en => width_counter_enable,
		q => wire_cntr3_q,
		sclr => width_counter_clear
	  );
	sd1 :  arriav_rublock
	  PORT MAP ( 
		captnupdt => rublock_captnupdt,
		clk => rublock_clock,
		rconfig => rublock_reconfig,
		regin => rublock_regin,
		regout => wire_sd1_regout,
		rsttimer => reset_timer,
		shiftnld => rublock_shiftnld
	  );

 END RTL; --arria5_reset_rmtupdt_t3m
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY arria5_reset IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		param		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		read_param		: IN STD_LOGIC ;
		reconfig		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		reset_timer		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_out		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END arria5_reset;


ARCHITECTURE RTL OF arria5_reset IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "altremote_update";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "check_app_pof=false;config_device_addr_width=32;intended_device_family=Arria V;in_data_width=32;operation_mode=REMOTE;out_data_width=32;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT arria5_reset_rmtupdt_t3m
	PORT (
			clock	: IN STD_LOGIC ;
			read_param	: IN STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			data_out	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			param	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig	: IN STD_LOGIC ;
			reset	: IN STD_LOGIC ;
			reset_timer	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	busy    <= sub_wire0;
	data_out    <= sub_wire1(31 DOWNTO 0);

	arria5_reset_rmtupdt_t3m_component : arria5_reset_rmtupdt_t3m
	PORT MAP (
		clock => clock,
		read_param => read_param,
		param => param,
		reconfig => reconfig,
		reset => reset,
		reset_timer => reset_timer,
		busy => sub_wire0,
		data_out => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria V"
-- Retrieval info: PRIVATE: SIM_INIT_PAGE_SELECT_COMBO STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT0_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT1_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT2_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT3_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT4_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_WATCHDOG_VALUE_EDIT STRING "1"
-- Retrieval info: PRIVATE: SUPPORT_WRITE_CHECK STRING "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WATCHDOG_ENABLE_CHECK STRING "0"
-- Retrieval info: CONSTANT: CHECK_APP_POF STRING "false"
-- Retrieval info: CONSTANT: CONFIG_DEVICE_ADDR_WIDTH NUMERIC "32"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria V"
-- Retrieval info: CONSTANT: IN_DATA_WIDTH NUMERIC "32"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "REMOTE"
-- Retrieval info: CONSTANT: OUT_DATA_WIDTH NUMERIC "32"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data_out 0 0 32 0 OUTPUT NODEFVAL "data_out[31..0]"
-- Retrieval info: USED_PORT: param 0 0 3 0 INPUT NODEFVAL "param[2..0]"
-- Retrieval info: USED_PORT: read_param 0 0 0 0 INPUT NODEFVAL "read_param"
-- Retrieval info: USED_PORT: reconfig 0 0 0 0 INPUT NODEFVAL "reconfig"
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: USED_PORT: reset_timer 0 0 0 0 INPUT NODEFVAL "reset_timer"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @param 0 0 3 0 param 0 0 3 0
-- Retrieval info: CONNECT: @read_param 0 0 0 0 read_param 0 0 0 0
-- Retrieval info: CONNECT: @reconfig 0 0 0 0 reconfig 0 0 0 0
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: CONNECT: @reset_timer 0 0 0 0 reset_timer 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: data_out 0 0 32 0 @data_out 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria5_reset.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria5_reset.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria5_reset.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria5_reset.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria5_reset_inst.vhd TRUE
-- Retrieval info: LIB_FILE: arriav
-- Retrieval info: LIB_FILE: lpm
