// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:02 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o6Ju3v8betvVh8Wn00hP87VMhv2GuE8MNlAGiLmvV7zA7y1F3qD/EbrloIOCjL4a
bUEUNm8fx1j5ieQjBJB6lsficm/R3vSt9KZC9ssVxsqDZRNafk/ml/c9KVMrwQTn
k+VcWpt3GLyJeg3BogQekLZKUwRvQj/E+VMzkwPksdc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10528)
wpc9/HptrjjxvAg0FA7PD9XaSLyeeBH/I4bY3XmR3wLr5iXZlD58Aqq0b+JW+upu
W8VGXynCx7H5UpnZsFNzhyn5sc+b32QOahT/fueQ6imZ1VGHaMfresg6H0/GgQ/x
nJOx3oi5UDQIPV6bYMXjis1G/Px7eJDdZjO5iIbiJfvKEKXeHy4etJcTNlR2WuaW
Owc2bbt1B54RWTxn86pxiahS4cTw2IXghLA2FHTmYZeYK6/Jz7bkGA7zI755Dsvy
1lfzZtvVXGTMIs3D+WM7t084FFc/t8YejYOU5ua3hkqF2IqSVsXY9F+ixMUc1apZ
KB+3WK+brm36d392lMzhuQsLfk9Kw8AnuzG0g8x91SV11yuhlzputi+KvWptsBU8
KSaWxx+z2b2eUaG677PxGClU6vY68g4uQb+0w1VMvkbr/t+4q+9DH7ydJL2+XmUG
7dKGtdB3JduTjP6uHa0ClNPAM32BqveR0+omGqR9UfTMNQCRm62MrRhtax/bCMCy
bz2OgAlnrQ5X/bhcdhI9QX8pqsOukUigEupUnAb0NydiWzUQg8DHE9PT+DK1v2G1
BXIvO2VkuVmNh4TCQvFqp/SJkLUIbZMd9AmeSxYtheeuW2VkZHSEXR0U6jkgDRfd
J8aVO/PZ2Esx9lGkhLtPArAMio2yedf2lEtM29yxW1y7+eh4BESN8ofyPTmMwsVr
QNaf3Kp+NaNLhzQf328WnGYGvjp9KiEa2JKmEyV2lahCxvVX9TSnZS9eFxtAa78O
3lstWk6rQOyGW99x2mMagPX8/kZ1BI6uZiUoDO1s5rOtXk90rOcDRYcXCvZHe16b
dTS3j81JU4ekU5m+A/JYrANkmGN2rEOLu/mMUWSF+oWRqQyHiSWmtgGNXa6PCXzS
hcscMRANL5RpRsF+hou1rnnMeDwGmdSn04OI4KHuqooOK8W13SAu/lbt+GmI3YOf
W2LTHHWL4xs8khu8POSlqLIG4zM6vvIfAIPWfEYxsUKR9L654RQlrIQaJYYrKFQL
sPEnmMWVGdYoWfKHp1ERU1ldFT3RiwtpkSu2A0K080ICal/uNtjsCiqLLlRzQQbe
dB2398wm4uEQugY2BQ23MCQw80jEcCRBSY2a0nM8lhHyY150UiFBeRiY0wHrYikX
jGGJ3UDhumIKUKCYmpYhrPTHhsaYMSKuEW/SD//swtTK3LE5XK30metSJzxLKvgb
biBZBJLECx7/GSN8DQi3OAlU/LLIB3wRe3DPseF+kS29SNWJuXqm07tRSFHRgB2I
9kwaSL+YjMAR3iBOsqizONgebZ9KKEO9fqu2teMunh6LvbXLzUHsy8im5wQi0zC+
z/T/WFCeOgsZoZxosZ4LwA8Jg5LzwLtGFEIW9jsh9SSyD+B9kA8G95wv5ehlidIE
Bl0U120hq6bM5ZbGUI4P+xbvo1bFGDDFOEE37KqjRrPjqyjWFghK9wQ4RS9LrVfS
I8BqlYl+goZEdNMPTUtNCxcbXrSZzG8tGBs5ajcNMPHqWsFCwiGF5/icfDhP6ZPC
eEwQvwBFcDhmjM/unu0Bl5wb5EfXvMFRrGnE2ol8BaOzL8glQlxV8QraJghi6ATs
qjBpkdM526jWducyM5oPWkShXIHnS/0Cf7OisqiNe+C4CUB17XWYz4bPRk1Xg1EN
DoOsaIkXSeIO9LZWsCiUQ1K3FN9G+huZqLxiwvwGBRA0bE07zODwEDNIrixfMzEP
s2hwmdFnASjVJ96BoxbTePhJ0WL5YBEj3Xh5WOBPE38xbqh/3dZ0bH9d9d2wD+wR
7WVU5ZxCRhK9BcZR0TteE3aHVIUiTQ0wCe+k451mV7dtW96qaOFaAHhcBfoE2DcJ
HZYSrSQ089Gt/w5N0gvZy2oLUkbIIBh2lXnadUs4KZ1HdM3HbCubSNSf/LxHdXq4
C18zcvrRmln3FBHulpK+4YnX/Mk7Q0zErgauCodv9geXaeLCBiy5re9sJRhBJzXu
nBvypoEpkZwDY36F8Hf9xbsFKyAWGgu3uW+geCtdQWRbd5ikdRLZOaNXocf9mKyD
G4HmyRFCyNK5djdD6iEdA3dyQhWw7bS9SIjZeR7jtQ8E155pbX7PipCH4HZD4Eqa
vRieMeaSl739G5fRA3R/tJOsVBlbLFVH7BN3CtyEqHznFiXaO25/k5dT/Xl1Mq/U
VeG/t5brun78KlSlYCJEQtgQhESw7M1j7BDhmwGrCuTaNztkvXqbQpximpg1CgyY
TmA+nlnsQCpXH/185gnYq0J3Q2OuosJVocoVIMaIENOz+ivNI0LgaUEdUdUWd1f6
eF63CTwZG7ggMGJOEyUoP+lA4weNGvwb4Kcs2aTbRbl10UJCZ4l6geXngWknAGL3
Pa+4f2QcCINWMng0LwFx7Mhrm7//gYJ04uAHx/kCDaAHLPg+4seXLrTWmHEOa1C1
CdB6DUNHhEJP9S88lIu4j+Q9/9DF80a+kBgqU553LaAN9Zb6mjIixAZ5HwRcn3wX
J93KgbxSMx3sB1TSbS0jhHaY6ueyjwHanPf2BKDvuLnpuXL92sExmKifm5zPGt5v
SHaGyTpt0sHGo1odJwIF48QCF6ElbIKooVb+LYvoueaIZMJmRYIVyKCfVIx6Jm9C
WsbAccTdChwzaRc7V+A1vfY/wolF84B3lBH2JyyIWXYDm0BKMvjUKmU4+zcS8BYo
DwwWBaDiuxIMpNl6J7zEQPIsexvciQqwVf/UUpvZ28V6NyONTuMNhIxbctyjhKXE
0W8z1xGHjEAQX7QsXdIIovs/2fSG9u7ou/igzKFSkG4BU3ISp2ijahJEool6Mqsv
25CF0TBho+hvqsKXQy+ecvdsdJHmX0na/mlE30OjqXg3Zj/SoWT8bsqJVa1vDvBV
Zyl7clMUgadrPlam3KaQgS7tAgm4xDnOwakvAOKM5Py/3VK5Arlzv9hJJRT0YwlR
5BZFG2dzZaiTaE2qNU7Y3U5geY7TCVBs0IkPbz2Zk7zEP6R6avdaLOup0OQxuPRA
hSqg5nKr5zlUDkhKptFdd680ih8bnIvXuYgFNCSSJx+jPxF7vQ6kuPXOKz9RLp5X
6BeBhHw1x3MB0jfkMrqwtI0Z1e4a2AwgQy6HEC5QazZRZF6qMITun7fWzqypgQU0
tiNOibMqC4QipvjxWPKOYSLSE4u2Ja1qGDeDfaLt5LTPnvFiaQe04i2pebdKqOoj
WI98m9e7VqmmEwxGGEDbe84kcFR7abppJbVepNGYFiS+zamGuvWS9T/JVD7y/jP+
Yll+A5UgMavURC7f3YUiTFnPqUch6YRcftrLs8N8ooyoqzegww0MTrpAPgHbO7vV
eaz8lca53Ai0+w/JclBORC3MEdiLZXUZ1OrnCbqc92QmuTmrqXvrq0OzBspMktuO
X+b8/nc6neIdeW0rXWeMWWYjxveiGUQ20JGA6mK/B8PCTzeT9vfcFVyGLcTCI3HP
Ms12xfLh0xEO+Ic+nryaINBJLgAyPYKOBqDQGXot3HlkllZl4pV0iqW50mPGxSve
Pl0xVK5OFhCFMs9u3bu5pHOad2J2LV7N4eubIFC3cS3KgYnGEQs4IrfD7sSiXxVR
rJU0Qu1uAAdvTB57091E17PUJm9kl6eV9irH2SnXTREnkJORqoQPwZzLlZfeTAEb
5LGJb6gPwLRifXY3cL1AvYZ0UVsG4NipMmZ4g7cwtE0HcfXHx3DgSWxg+XDQlmOc
f+0oS4JmyQeBOCH1WIkmy+LVg55KxqD5BmsQTnz0gfXy2XV+c3qkcQBEnu/3RZn8
uJin9C82ZccdjoNZRpGTm+87ucQhmdMAs8KgncxaGsbeNArKa1aMkZrWPkIbReZz
rm3NVgqPe1zYBf+QdlDlz2mQ/KO2rKzfmbFC5wKE3lQS7y2xLFCa9aPDbXadZOVt
WCuSdse0DbpLZqMN1wTmvWuqfMTcZLeWzEuW0uchjBXHIlDsfkCra4VNEn6qfbRm
sxUKvHDeni+pBmKRmASgGL/7SvaT1Z574FDyO4MtQQtWhCj6QpHKZsD98Bmb6gtm
5kNB6OkTbmcyh7fEdR/Zdl2Xi+orC++TBJ6n8O6nEo0UxMHMvYTb5C423Pip7zL/
vWilIyVJOj1WnhWS90x3wN1mHFox52L5ELJVBa2Mv2GaEdam59M9+wQcj7SXB1H8
1HKuQp6W9UQgwU3gOZ9jfk30OCyRSdoMznmLD8AzL9aTag9LPwuhWf8UhqM+7QvM
8qJIxHlx+aU2LMt/lvPfZru2+i+0qVCqIr/spqxxBpBkK4f5/OpE5vRL1sa5+C3+
WczHhKii2Gi2cX1F5wxye2uVp0rRuSVYA1M3N35hGLwLrkXV0LlHpoq51YLoB92S
avVYpbrx7GoTAILhKF8LdNf5IlGcMXRUWXpzCAHN3/YDHhw59iROzicEvIHhcNNv
vNL4xQ2P74OJ+ohWnlB2rt+lH1yNgvHfvPvb3tZzKidevF3tmnGL3nbGqgqkU7FW
0K9Fffyg95Cmco8nhFR06ECbgvw3PnrKo+4LdoIzofc8NmeL0sPpGEG5l79jbd76
5OGKJjxclKRPYtXSE21am0Sm87BQ6jSHdot5oxrRoWRoHFr4UrjL0cIYZlWxyoQP
5WdNaCpQYbN4JPXHk5RB4/VmqmjHEM/WM5JRgfLhq2hW6N7SeaHcFTt6A40Eb3Es
kQIDZUbUSBZ3fk+Lkw1eY5dAcWWrC5Zvnkp4SVg04/+/CSrfpiaQJWHlKN7gMG79
uyYr5/PVDyAKiECtOJNslZ2dLVKbNNCHssGtrv59MYNUyxTJJZeab2TsP8whqhDZ
ApsQi6eFTYOYEVdVoFpeP/s0icmOyF5AGgnam8F1CYu1wWSRONPPoToiD4k3ns4O
RdC24lVvIrQa/mIMZsQvbW+M4UUV/muA5dvaN+7bbhnnG+ODsfOLqG/9H8c2W9No
alMzGB2CncGLZFMAsHT5d5KDpBr8GncfHuZq8RbGZA92+h11ZFp4OCoWXy/cPs28
UE/eUFgDi92adQ0JR3HBX0id2jNzXwTcHzepCj4t6TKkAK8/acsO6kIOWLRdkI1/
+F6wgUHOH8uj9gXYA8UkKBEJsPetmhSISvjoXtcNZqd38sy5Uuqu3OrHr4/tYhG0
3rSSE5EXxfs9HorfY68CyPY/Uo/S5qc1LUHrB5lzPiS0EkqZJtlCsg09KdSC77SB
keDNYGDlJUqvEsxVAhCS3OjAfgnU0c8chufKObBIvxGBkRPq98nTuzi6L4tTHYxn
tF8gX1T23t4Q5V/P5YECChtuogdwAJZO8I4CqVnPgBrqx8PtPMJdqmG83fmsY9gK
6o97DBjTz1Rfrs+j4vazESswlHkf8NdjwXwhy7z3ZAd+GU7UhPH3leDjvpmJ1bfD
aN6Wtz1M6F2p4HitmxGnCAloL33cosqMZchYqhQ1X4cCLZTLnKC2OBJxaIvar1ok
9CrWKF47LnKyrfPXEYs1m0r1ToK4nOTwHbWzIsrsaYp3cCPnbWtn8+2aAVIGAnqg
RXMiVwT6h2C1QalxUPHCai7sGRdat0yXrvWHSTa5q+uMCYf9zXmjAb4SR6MRTmk1
u8YnwGgzJRmqeYN501s+ttUAeV+9NNfXuJQePvihKhVhaTuPS3thxENZBGL1SCAf
2kyU+3wJ+adXhA3r1DD0s+yaxVGHgL88oOf7mCaRUrrva006AlJuLvIpAEisMJhP
e7rJwH8N2daPbleIXbQN5ltppwa7ilGL2TVfBb0WtBEGfOqw/qKIsalURuFmAe4I
WAnNBtCwSdAwIMj4gtwim0YTsCCmVFr5+yXCtqCnNfzjRotOCqf2i5/g0MpHMsZE
0z5MNvMsqJxR0RSXLjkmN6hdttItjwASgrNuRGr6r8dNFEjnLnFreKQCne5sgb7r
oDEFZAyKkiIuCw9ufjcT0lNKtUBVC6DoYi9cGKlBdpF43WBTsok19KKPmUjqOCYW
g60DMLIhR0lng4NQHExTJEGqcbNzhlgnGQz0sEVS5FQPUOjtP77L0frq/VkU/++G
4eWp2HOkz3sNTNf/8A8WE77zMjxPp9VPeAJPGZBXHPFwlWRrExzwCk0enEEEXyzW
Pv6vbrKzrxi4A8CDJqboYZhFSnn/3B/OXEb3pbpabSx1niA18trj5H2kg1UamAdS
FQVxuNNPwlLcxABeavGi1BBaVlNwVOzACQh1mlukEjDOQwSP+ZlY8YfoPxdbwGRU
rQW/tT+rQ0RumB5Q14m1CmAlCTuH+zIBXspmdGHkRsVT1gqm4KVjBJtYesHhSsqN
7CxUkfkWd5W26Cb+rP8T63NAZaGgEtXU9oooaOdlRTc9I8k0QfrRfUo+aEsli/7p
Eum+saPhWeQzIzu3scqET4UIDzKGnb4JRUZ7U201CprtAbRMb8bT+iUYNxMebFbn
X6omzvzWLmz7Rxz2jvUKMpITsE6u3GZP8yhfxmF1xNpRA1fwA2jnrIDTOdMiAyxb
/Wo8swvdkXuKXtHqzw4FZ/UFHbQH58E5ucDydMA9v1mloNhZhb6hXTWjTbF1Dtc2
4xaM5Nc8BTpkE6e/l6ReLvOz+w3YUWkb+SrwqajPBYN2sYJqJAmvDcHupfII/5Ps
lXvzAAg5ac2PiPDPIisu7alyAHFpBr9vjx0nMpc/YE9AeVdH+zh2qzV/q6xomn+Z
b4tPmHlF+Fv/lKlMDcVfP+j9LD2tpl7RWoHl4ItVYLTwyX0V0res/3jyc4juz48/
b5lane3DLYbQU6uiVf1HDGwnrE3njcmPJ33uRPNPBgMbzV5AcZCQc7M5GxzQeeHe
lv68sBhoWCDojoxHtSWbXsiNjzatRNLA+H/Nnzc8EfYwjv/W46k/Alk45s4Qjzqn
85l3fmAkokqdATsVeKJ8nVv4Bkt/vJPQVT1DUgPZqDkksJhitZJ8olsbEs4z12e5
XKxAR7nWPc9SIddEus9w57DVJhnPQd3qD7tTUKE0qfM+H6Z8SBx3vypePGR8014w
msA/9MFdHJMyhRVDEkNGdJvhK21CHekfaoUnZv/xzJK2RVDkQG/yo/yFIvZjAb/S
Y9/QF+D96gN6AS5Jo6feMUB/6NxFqJqo02GM4apONIHbHJs8gD8wbDg6r2hBR+Ie
gdGr5GwpmJwBLZy/f2QEXWxJHMBXejuhUM52MWCj6H+4022xD1L79l2SE8WpEyNU
0tVr/EKiquwTheGAin/y7XSGQn61n8DF6lh5qEwqlttkYYVEbUZlrbEX+jCNzjME
VXtQ6fbv8dLjk3XEI5bCmZwEnpk3/f5y4f5ljtvL9CSb+/ptdeD5c/OyBNWi+IYr
u1IqoqeJYm5kn2IkeSEBebE6IWCeOpqIjwzjWd0OxTOpQ8iFVZ1JhbbSF1U3DAvY
2zRT15Ura1YeXqtwbX9+s2Cd6v5vzVCBRoUWZRmxPjeN4sDWMYzf4z63KHCOjPEF
ASgIEeYF4L25iQzyyqXMtbxHpih91OwiQKJk7sd0UorbWqfyh+vRQKH8+QgDBNXo
/Q87rvW7Yyr0FJVldoyqQ365xcMA5nNKp3mZ/ToJdo0tPjiS4YcHtJsjX62W8Cds
m5qS5RYH17UpHQX1RFY/UzrxuPHz6Yd5b9kGAb3+keYrVal3sMuYX16U4lq2xno1
1ihJ7mzvYlR9BvTNp0jbfthpn4SPOvsWhfHcEhkZaU7uNyJRjz3QfpM/7+/QQ7lW
zvT3B/w7Dn2ae0ZgUTjRWZqNuoXshkZjjsRE0WRolgCfYA7uUc1XPmq5kuuujZL/
AoypXgM78FMw0j8J9hhwa3DHhiYmDgBJoYc+ZaOcS8snuAWPKcpFwID85AXK1jWZ
baOd5ZluWtyAF26SOgkuUFVIti5c7ynIGIst0S7TZc2N1kGtzDOxT++ME5rtQB/J
p8ltw4STDhvVz0aEeiNkZYD6WnLJ6ItcbzhYoa6KkLbtcRZn6uFHTQM2A/HySc7Z
EGp09UNIY3UEfQiY31fNLiK+bpy7MV75PVMr5SjZXvZVGV/5UnPKl4rZElnFiB0Z
JPmAcGkUv3gLsTxHUg4Gp8hQ6MiBpbIp4x0IMkd/OtPNWAz3i+qj+Gwu2gW4cPxM
5XZ04RbjV2I0WjqWYU8iDHPnFwYp1nmCXQhCI8xjuxM4TMV5iRKkqFGY0mhpFR6/
QBf/xN3Gyt6NByv6Tb1AXZc7ppohtiGNAouxa+IfUtEQySaGSwDkBOA9b0zKxbGq
cOelK/DfC9H344CHvGkzVOI/vKBxDXIg9dAqkxQ3AtP/2DqjY346FCNnmEPkC61L
VISCJmRTj8+mUPveztch2MamwZY4n/bOhOkuqKbyGlkLtSq/Vvu5R45BsJEWPXqE
Q4A9gyI2ELaGwRShJqjyE714gd233xIwaxb77p8D4ZSMKU4brQDZyszoV4e74T5U
zhBWEjkzqlJuso7HFfQ2jAavgUZCvQyLNF8VrvcXn/mB5YY55r83ZuDKH78E45i+
nsT0eupNrGahaJDTY9n7df05GVMifEPyO5YnrvkQ0Sb3LHtWPkNMCDYnGr1QDfb1
TkzkIXxj3nqZdHmiWYhJUaZY4xgCaG31kdOWSqK1yVFu6wuwMWgOdOwF4h+KaIIx
hpgr2fzkIjfosKO6+ez8CbU6VVo8mwvmHIBc2bHNoxoKi4fkKLEq4xiURVmxsaiD
voCUQemCQ/ibZK5IP10JTW3XN11MCLdJKTDgD/26NeP5iN9xAwOuKE70y52SEdez
rp6lUZfZL+P76UdRMI1PRL0G48x+xb6RNV7149hyMA3H1s8HuOwhFHZwiUadC0SL
JNyk36MDAD53e734Lb8Y3CbrLqdqhRes05XRzPx2TnzSGEx/irw0CQAXmiWdXK/h
qKHC+pyuYNtnM1fBpbeFUX5XxQl5/QHEZ1pGFBJ7qLu0yZcHfr3mxFl1EN7b2Vo2
DIGHi9b9NhOqf4JYZjD10q320JAWh38LjnrM5WUu3kBM+s6GvSrB36f9lAMnzfeu
WZ4+zQy+MQ9LZV0giL19Nuv9T/MvPvkCu80q4hVwsTUoamnEk0Mck1nSNUAX7sNX
uG6kywY9hpswj7fp8Bw3KhFYsn05lbER+ibJgCvVctyHvuSEdR5g8e9ZRupJVJeS
G/Bj7RuSgPK6HNRsV3B14sTgSoOfVBfuvp1pE9VEKAGa9n2mdfXqFVyvU64RQWzv
nBlh34QkghqqgIEHbVZDDWhjJ127LcSH76GcdfwJINrUX0YW+vYrsbHPdn3Dit0T
+1FY9eI37rVTkyG9DxS2/gOcb1CUNwXJDWClPCbkYQWXsRRUZY71B0iinNWv0Sb2
Vm7RGKKjHsBKlyGfcAgOoio36VLxj/LNZTUGH+pv3rhpLHdoxo+C5oJqq5MXKi5k
PXnYUzbgsRL/aDJ1imI7IeX1Zdzm4VlZHNz/xD5ccnnvqaK4Q5pudW71HHBs44ee
73VRbLG33un7Sl6BnyrCdSGApcAvOoRg4Op1huax2ur1dnYvB6VImWkNGy9U0fM4
GT97UMxpJoSCym04uUsARGIyHkMVzn9SAZMvvD6Ub7qV/1M31iculYIrDBF6sIgK
vuLVygT8V55N5PmEXTPGzZki17ZgFq4Oajk1Makms6elo17xE+9nv7yKdiEbEVc/
3pJumydDxT3hiWdF4FRYKHys/IJAh0nUK+Voyfybtup3c9K+u3MyOK1wnN6jJyrT
xds8kZYtWcGOAY9k13JDcNp0+4Hd0yuyWBOuUTKTt/LIXSrQpXapPmGbkMZyGMrC
UfUJtiTmJC6pbLO/pih+tvTE3RCDp4e87shR2gQhDxDbtNZGpH4JZGe9nG9RvwSq
6TMbI+DCCub4TPSudrzqZaB89hcqJ2bg8WT0ZorOpWTtODZbK0uwcatbClR/kIbx
uaD0jcVFY9tl5XJkjPTgjDXbNr/gXiI/mo/I3zkmb0JEqDVD/Li7tJVpKoQXimek
PHHE5j5hQh90P923hIhEjQPaydB0Qano5RZ2ueqnMrYRqnvmGRzHLTbEJC5LP/Aj
YPmehBcx1vbib2qA1xuD/EztSF5a0mjgXO4s6fph9I7JkqK+JoVcLrCISbwnyxQB
tVydgtqXTQme752bti2EziwbOG15bR6TO59X+CsLcJT9G1ARqj9PQZNE9NmKVoEl
eDT3bAZs3kG5gaRmQfoWs/N7vFlvezYLzVYCScrYDKZMEz+ASh641eeZhIq/Zdll
L3FAoDYDw/HYRk3dT0TRn5pa5xLLzFY0ylXgSviEgezUo4YgBRzlUxv1wlUbZy4H
dA0DHvRk+8DqoNep45Tu4XaWEk9bvuZJQRVw+ftMs0/OyLGZ+UW8dXHLITxmrEqF
IRlO4VnA/Vlek9PlXMWI6VuNG+aTWmxUR3U1Za/DbE6/5Tul7mJ7MvPL2+qEpw8Y
RhGHIJskkBNPqXR2sJbcj8rD67bT6jlTPB1No4H7Ux9v9VHI2nQw2ItHzL73RbAf
giBZnRCbesB1+DFVKciLuiYx5RdXxJ8qbIq12tlC8RZVd5y3fsCNETIjo5hKW9LT
6/D9/SfX4LeOziMxE5GPawVWwsN327kRG70DYN4QQOVMz90geeeJjH+A2l0XXpS6
C4DDbLveC5FtLsyDkDdIHTstT2jnvOATncnR5cF9mGlOAZBaOh2jxZMuvAxY82lc
G7AO1E0XB9Agz7Oi+hXI0TXzuYOtLOK9nMtP6sGYLZTqoj/Gs3vMrUhBAm0vQNNv
PbGiWiKb3BZ1HrnIXPHm9yesMNfvs8rZr7Guzp+d0i7beE0MgOFG9O3e37C+xxJ6
HpByWDIdXtTZrJ+YEW5+YRsE9B/e3oqKW46sE9FpTkn/lrhOFl2faMhl860Psro4
gV3RrWOs1gISsfjzyW4fR/wipSPe9ZBHIotKiNYm4fMdji4qstPB8qabxJgj7ua/
vMiciLAtlMx6W3Akk5NqbbyuPi8GybAoM99qkWdICHqoP7Fe7fDQdlluxuEs3DRL
myhzBUkcSSdMCgh718+IoS1K+TlbJ6h0mltL09gptd1zSXKlZKtn6zQ8XKaUpLbh
7JN1/8AzYTN7FrB4nisNsC7Yze9xrdLc0323ETSu+/PpmsW63BSwAMYyoZC9PxVU
R0AYeWrTF7i88rEGTMvIxFBCB4vZEXzW95LCvS13/O2WS4RdvSX1uFuNbHJ6CmAD
iuq4twW2ZLvAlse6y9eA/bCk7CBiQEq4C7BZe6dmf7R5hc38lu6K6HuLGG/RuJvh
iQn+BhF2nYTBxsZRNWgJNl6++o4Wu6W07Ow+uTwwS29uaOhdPY8p878JN6ez3BmU
tbzqCUZ+r47g4FZsYtT71L/PH23yi8TQVQAZXVz8SMIKeqLWcRENv6UQafDF/r/d
gwz9pVZ0slqBZnykOAqlmiRP3nicJyYxlEBlWE6L0y2DXp1qSeuqO3GHLRDpAC6q
DWZc44nuLmfPi22034zLJ/xEKuWnhJ+ghiJQVrEhyUHBEI/Q0ISXufTV9SRjnMNj
mTdhkXJxKkeIe4d/BHh20nxEvfdflCfrTvJK7ReLPTmAxE4kNY253kFl27meAN1Z
WGCUM9FeCAp1enykLseKAye3aebmEWQsPtfaQelkXYa5QtiK8UmCclyvrQQ/DVHR
KUY7B0vNoZZpUcRYCdqsIQH+qgLVv/Vjx/gWwV7RHY2jtPjclJGeyg+GfZFt3j7f
IWv81KJR4hRzITL5iGoBCxhpX63OzYIYLyJ0tp3XY+JE2PwK2ORIBaYFMotpM7qs
G6HJF2tZITxqlthqpGqdjqWGpkFpML+l6aePxVNcAFMhQQwGFMuYHnsD9G3rUoNc
8jx4S6I8OkyZwny18rwKGmaM0sfbBO900+i2OdQwII0bcqiLbSThTP1vDqJoCjL+
8JH7jffls88/QMRBpWOM79aqdUNMJo3MxTIFrP2M3tFBSRqOZGAgQcBP5+era1Mo
9H1Upt0RanWihoRcwAkhxLwl94O/PZsu936GPX5kpaKY4NZ3GbcWboubHANd1o/o
nbMLo7aYfNKtN0SAaaf8LusSWCGZsdCF7JmEdCcmjQOrWcAPne2kTTm9cXYAX/mw
6Vv5xFsQuQwj3FAs2Dj7jejKYzGsjFIhIl9HT6ZQF9k4xC9g9elHVaQQ9D6Hu79T
xV0tZbjOVxggmp1pLPVlOKlX748TBQ5ebBph3njwI/bqU3BRWg0NzcQfegQ+1dy4
CbfeglIQRGzzzU0yG7pFn5b/TTB/3iqyqB4Oqzs4q5+YCKxt2yFMHJHZqDwBK1xv
U227R2Y//t92883O+Hyc13VmioPRBf8w/PIHaO722vSzccPmnRn3q+LuArkV8xiU
+XkNQj2y3Tl6dAJn+JoJQZiXYuknR5LIBd31KbIM4AzmcLyXVnpwPr8KFp2PF210
u/7iqmOKYyJNP2xbyKCaCBcYc0A4jrxvkoCo3Y6ZrfT5MlFgsGwkR5ec58c77Hxw
QsGyrqwHAe2S9+8X9/BmFu0czU33JyMnwhMWhxzYT6kqSdd7KDnWS4kzD+w5df6E
SbszOwy+ldC+Hu0n4PiIrlb7F8qvdvEVpbeqDfOyFoo4M6NKOylXNRWgoCvwEWaw
Zm1q8oVCo7RNuoFUcIQsexMYJY+U5/szoQoPYRQJrnbQXiVvaX2D98UcWo0Pn7J2
sXZTR4bD4fuul0UFgDAcGHWo6dS3Q7v/HS4a4jBwkWTSgs8a7VloT8qCxxDEJ33N
OTgduV2Or/z3GIsca3BpWkhe+AdzbAvnXeMicIK9X76uXSb7l1II/pe1QcM6zHXf
2RtS+QLDxm296jihEzKJ6tr4IZH/uC03Axjo6cP++ZZtmEpcx0Zxh/1syr7Coxx9
g6ziXKG+to/OmgBcPB3Zvkbueenf1/X5w76TzNw6GvoYZGDDcbiZijIqtv++vcEB
TKfq5KAG1ko4qb/uui6A5XGPvl0oqsHit8GVjUTI08A4GfBp6nBW+bN1jV7IXWGi
ZS5cs2rhxXMuUDaJKmresCskSy/L+KTLmICq4o6PbH1OB94/6T89EUizf5v7cJe/
4fPEeVDoJJ0VT8/WV/AnIOJ2V1F18wjoJurTtrHCkv+nUSMmzTmA4RFP8y5Ev4RX
XZ5yB89G/aiBx2LPq0KvuE2vKiOdhvnBiWpt7hzVWt+QEu7jnSSzZ8gvNDYwbT29
/u4xK5WltptnuFtvZAz16vcRDcbFoZSmjMm4HgMxkPTOgzRfEiVTMAyvrhUS0g5n
zYN4UgHbQePvc09daU8tYhmCszuPPwfZLtS+GC/zdGeQObnZBQo9MC0Y4CrXayQa
3azzCIPbaZ0KW6pmmRuLYnWhxPCV5+5BWjHnxRfzWX0S0y48crRgnYzC/CrHgo+x
sUlne8AIBBazLBlKkKEdam41A3ydVBkNqysL4j8vUYGhZif535qi4w8fFbH2oITM
WovU4xg0pi0VyAZtRDHilk9zDsv+YoaRil7IODS1rPPVva4VHY1COgDzBgM5eQBt
oEu6QxmwPGzLrgjfCReN5OBdBc38l/U+5h/Yfcuyx4kZ1Be3MMoqsid6L1HXkP8j
ngT4PoE7yJelxTheOIZaD6RRs1g0L3M6oVDHuIRGj1yYFEeuGrNP+RbihF/TWdOC
i3kzS52Tn2QvQFz/M8PQneR/ZEd3PLJG111oxe6aNY4W5cOrk15VLtuxsOqIEu8n
9/P8ReKU3JDvwR2eSKjCGY5tx3zSVIH8rPfT8UjyY9czYtJUpjk6I32L8xHRZr/r
hy0cNqehKnz7FOmzI3pZFRQDgQ1/h+1/gacV1iKlGzot4WSzuWgZon80t5fUBuJ0
XTtyYiHcRqP3suR5OKF+gXT6iAeNcslbGi2ZX1nFsafFPSefEUubmG/lVEdaEzOw
aKIDFXmqXCmYg+sL1dNxHYUdTFozUxOg/xrIUablHNKWCAk/Zj48Cu/R4KYDZcok
UnOedQjKrPATfEJsN6JHD0WVlw7ffPkHquWVPj0r/D2777tW8nyNWl8VfAi48Gil
jbnvU5BY2Nag10obqA0kXRrH99jVm1Iw2y5fd7DBrQ5fbrjnZtxYXSGckpnOdw6j
iNLgwK8+fwF6+3qIWCEE4g==
`pragma protect end_protected
