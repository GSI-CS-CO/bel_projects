-- temp_sens.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity temp_sens is
	port (
		ce         : in  std_logic                    := '0'; --         ce.ce
		clk        : in  std_logic                    := '0'; --        clk.clk
		clr        : in  std_logic                    := '0'; --        clr.reset
		tsdcaldone : out std_logic;                           -- tsdcaldone.tsdcaldone
		tsdcalo    : out std_logic_vector(7 downto 0)         --    tsdcalo.tsdcalo
	);
end entity temp_sens;

architecture rtl of temp_sens is
	component temp_sens_temp_sense_0 is
		port (
			clk        : in  std_logic                    := 'X'; -- clk
			tsdcalo    : out std_logic_vector(7 downto 0);        -- tsdcalo
			tsdcaldone : out std_logic;                           -- tsdcaldone
			ce         : in  std_logic                    := 'X'; -- ce
			clr        : in  std_logic                    := 'X'  -- reset
		);
	end component temp_sens_temp_sense_0;

begin

	temp_sense_0 : component temp_sens_temp_sense_0
		port map (
			clk        => clk,        --        clk.clk
			tsdcalo    => tsdcalo,    --    tsdcalo.tsdcalo
			tsdcaldone => tsdcaldone, -- tsdcaldone.tsdcaldone
			ce         => ce,         --         ce.ce
			clr        => clr         --        clr.reset
		);

end architecture rtl; -- of temp_sens
