-- megafunction wizard: %ALTREMOTE_UPDATE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altremote_update 

-- ============================================================
-- File Name: remote_update.vhd
-- Megafunction Name(s):
-- 			altremote_update
--
-- Simulation Library Files(s):
-- 			arriaii;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altremote_update CBX_AUTO_BLACKBOX="ALL" check_app_pof="false" config_device_addr_width=24 DEVICE_FAMILY="Arria II GX" in_data_width=24 operation_mode="remote" out_data_width=24 busy clock data_in data_out param read_param reconfig reset reset_timer write_param
--VERSION_BEGIN 13.1 cbx_altremote_update 2013:10:17:04:07:49:SJ cbx_cycloneii 2013:10:17:04:07:49:SJ cbx_lpm_add_sub 2013:10:17:04:07:49:SJ cbx_lpm_compare 2013:10:17:04:07:49:SJ cbx_lpm_counter 2013:10:17:04:07:49:SJ cbx_lpm_decode 2013:10:17:04:07:49:SJ cbx_lpm_shiftreg 2013:10:17:04:07:49:SJ cbx_mgl 2013:10:17:04:34:36:SJ cbx_stratix 2013:10:17:04:07:49:SJ cbx_stratixii 2013:10:17:04:07:49:SJ  VERSION_END

 LIBRARY arriaii;
 USE arriaii.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = arriaii_rublock 1 lpm_counter 2 reg 43 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  remote_update_rmtupdt_6co IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 clock	:	IN  STD_LOGIC;
		 data_in	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0) := (OTHERS => '0');
		 data_out	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 param	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 read_param	:	IN  STD_LOGIC := '0';
		 reconfig	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC;
		 reset_timer	:	IN  STD_LOGIC := '0';
		 write_param	:	IN  STD_LOGIC := '0'
	 ); 
 END remote_update_rmtupdt_6co;

 ARCHITECTURE RTL OF remote_update_rmtupdt_6co IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "suppress_da_rule_internal=c104;suppress_da_rule_internal=C101;suppress_da_rule_internal=C103";

	 SIGNAL	 check_busy_dffe	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe4a	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := "000000000000000000000000"
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe4a_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dffe4a_w_q_range225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe6a	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe6a_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 idle_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 idle_write_wait	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_address_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_address_state_ena	:	STD_LOGIC;
	 SIGNAL	 read_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_init_counter_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_post_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_pre_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_init_counter_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_load_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_post_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_pre_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_wait_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cntr2_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cntr3_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_sd1_regout	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w431w434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w431w443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w437w438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_idle477w478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address179w226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable70w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rublock_regout_reg529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_range173w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range427w445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range427w440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_all_done505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_param_start_match485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_param476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_select_shift_nloop528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w8w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_all_done489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_param_width_match490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_load449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_param475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_wait448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_range171w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range427w428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range429w430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range432w433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_idle477w478w479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address181w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address232w233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address237w238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address242w243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address247w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address252w253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address257w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address262w263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address267w268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address272w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address277w278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address187w188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address282w283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address287w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address292w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address297w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address197w198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address202w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address207w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address212w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address217w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address222w223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address227w228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable67w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  bit_counter_all_done :	STD_LOGIC;
	 SIGNAL  bit_counter_clear :	STD_LOGIC;
	 SIGNAL  bit_counter_enable :	STD_LOGIC;
	 SIGNAL  bit_counter_param_start :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  bit_counter_param_start_match :	STD_LOGIC;
	 SIGNAL  idle :	STD_LOGIC;
	 SIGNAL  param_decoder_param_latch :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  param_decoder_select :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  power_up :	STD_LOGIC;
	 SIGNAL  read_address :	STD_LOGIC;
	 SIGNAL  read_data :	STD_LOGIC;
	 SIGNAL  read_init :	STD_LOGIC;
	 SIGNAL  read_init_counter :	STD_LOGIC;
	 SIGNAL  read_post :	STD_LOGIC;
	 SIGNAL  read_pre_data :	STD_LOGIC;
	 SIGNAL  rublock_captnupdt :	STD_LOGIC;
	 SIGNAL  rublock_clock :	STD_LOGIC;
	 SIGNAL  rublock_reconfig :	STD_LOGIC;
	 SIGNAL  rublock_reconfig_st :	STD_LOGIC;
	 SIGNAL  rublock_regin :	STD_LOGIC;
	 SIGNAL  rublock_regout :	STD_LOGIC;
	 SIGNAL  rublock_regout_reg :	STD_LOGIC;
	 SIGNAL  rublock_shiftnld :	STD_LOGIC;
	 SIGNAL  select_shift_nloop :	STD_LOGIC;
	 SIGNAL  shift_reg_clear :	STD_LOGIC;
	 SIGNAL  shift_reg_load_enable :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_in :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_out :	STD_LOGIC;
	 SIGNAL  shift_reg_shift_enable :	STD_LOGIC;
	 SIGNAL  start_bit_decoder_out :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  start_bit_decoder_param_select :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w22w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  w51w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w8w :	STD_LOGIC;
	 SIGNAL  width_counter_all_done :	STD_LOGIC;
	 SIGNAL  width_counter_clear :	STD_LOGIC;
	 SIGNAL  width_counter_enable :	STD_LOGIC;
	 SIGNAL  width_counter_param_width :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_counter_param_width_match :	STD_LOGIC;
	 SIGNAL  width_decoder_out :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_decoder_param_select :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  write_data :	STD_LOGIC;
	 SIGNAL  write_init :	STD_LOGIC;
	 SIGNAL  write_init_counter :	STD_LOGIC;
	 SIGNAL  write_load :	STD_LOGIC;
	 SIGNAL  write_post_data :	STD_LOGIC;
	 SIGNAL  write_pre_data :	STD_LOGIC;
	 SIGNAL  write_wait :	STD_LOGIC;
	 SIGNAL  wire_w_data_in_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  arriaii_rublock
	 PORT
	 ( 
		captnupdt	:	IN STD_LOGIC;
		clk	:	IN STD_LOGIC;
		rconfig	:	IN STD_LOGIC;
		regin	:	IN STD_LOGIC;
		regout	:	OUT STD_LOGIC;
		rsttimer	:	IN STD_LOGIC;
		shiftnld	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w431w434w(0) <= wire_w431w(0) AND wire_w_lg_w_param_decoder_param_latch_range432w433w(0);
	wire_w_lg_w431w443w(0) <= wire_w431w(0) AND wire_w_param_decoder_param_latch_range432w(0);
	wire_w_lg_w437w438w(0) <= wire_w437w(0) AND wire_w_lg_w_param_decoder_param_latch_range432w433w(0);
	wire_w_lg_w_lg_idle477w478w(0) <= wire_w_lg_idle477w(0) AND wire_w_lg_write_param475w(0);
	wire_w446w(0) <= wire_w_lg_w_param_decoder_param_latch_range427w445w(0) AND wire_w_param_decoder_param_latch_range432w(0);
	wire_w441w(0) <= wire_w_lg_w_param_decoder_param_latch_range427w440w(0) AND wire_w_lg_w_param_decoder_param_latch_range432w433w(0);
	wire_w_lg_w_lg_read_address179w180w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range178w(0);
	wire_w_lg_w_lg_read_address179w231w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range230w(0);
	wire_w_lg_w_lg_read_address179w236w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range235w(0);
	wire_w_lg_w_lg_read_address179w241w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range240w(0);
	wire_w_lg_w_lg_read_address179w246w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range245w(0);
	wire_w_lg_w_lg_read_address179w251w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range250w(0);
	wire_w_lg_w_lg_read_address179w256w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range255w(0);
	wire_w_lg_w_lg_read_address179w261w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range260w(0);
	wire_w_lg_w_lg_read_address179w266w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range265w(0);
	wire_w_lg_w_lg_read_address179w271w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range270w(0);
	wire_w_lg_w_lg_read_address179w276w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range275w(0);
	wire_w_lg_w_lg_read_address179w186w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range185w(0);
	wire_w_lg_w_lg_read_address179w281w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range280w(0);
	wire_w_lg_w_lg_read_address179w286w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range285w(0);
	wire_w_lg_w_lg_read_address179w291w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range290w(0);
	wire_w_lg_w_lg_read_address179w296w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range295w(0);
	wire_w_lg_w_lg_read_address179w191w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range190w(0);
	wire_w_lg_w_lg_read_address179w196w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range195w(0);
	wire_w_lg_w_lg_read_address179w201w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range200w(0);
	wire_w_lg_w_lg_read_address179w206w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range205w(0);
	wire_w_lg_w_lg_read_address179w211w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range210w(0);
	wire_w_lg_w_lg_read_address179w216w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range215w(0);
	wire_w_lg_w_lg_read_address179w221w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range220w(0);
	wire_w_lg_w_lg_read_address179w226w(0) <= wire_w_lg_read_address179w(0) AND wire_dffe4a_w_q_range225w(0);
	wire_w_lg_w_lg_shift_reg_load_enable70w75w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(1);
	wire_w_lg_w_lg_shift_reg_load_enable70w111w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(10);
	wire_w_lg_w_lg_shift_reg_load_enable70w115w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(11);
	wire_w_lg_w_lg_shift_reg_load_enable70w119w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(12);
	wire_w_lg_w_lg_shift_reg_load_enable70w123w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(13);
	wire_w_lg_w_lg_shift_reg_load_enable70w127w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(14);
	wire_w_lg_w_lg_shift_reg_load_enable70w131w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(15);
	wire_w_lg_w_lg_shift_reg_load_enable70w135w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(16);
	wire_w_lg_w_lg_shift_reg_load_enable70w139w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(17);
	wire_w_lg_w_lg_shift_reg_load_enable70w143w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(18);
	wire_w_lg_w_lg_shift_reg_load_enable70w147w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(19);
	wire_w_lg_w_lg_shift_reg_load_enable70w79w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(2);
	wire_w_lg_w_lg_shift_reg_load_enable70w151w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(20);
	wire_w_lg_w_lg_shift_reg_load_enable70w155w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(21);
	wire_w_lg_w_lg_shift_reg_load_enable70w159w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(22);
	wire_w_lg_w_lg_shift_reg_load_enable70w163w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(23);
	wire_w_lg_w_lg_shift_reg_load_enable70w83w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(3);
	wire_w_lg_w_lg_shift_reg_load_enable70w87w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(4);
	wire_w_lg_w_lg_shift_reg_load_enable70w91w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(5);
	wire_w_lg_w_lg_shift_reg_load_enable70w95w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(6);
	wire_w_lg_w_lg_shift_reg_load_enable70w99w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(7);
	wire_w_lg_w_lg_shift_reg_load_enable70w103w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(8);
	wire_w_lg_w_lg_shift_reg_load_enable70w107w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND dffe4a(9);
	wire_w_lg_w_lg_shift_reg_load_enable70w71w(0) <= wire_w_lg_shift_reg_load_enable70w(0) AND shift_reg_serial_in;
	wire_w431w(0) <= wire_w_lg_w_param_decoder_param_latch_range427w428w(0) AND wire_w_lg_w_param_decoder_param_latch_range429w430w(0);
	wire_w437w(0) <= wire_w_lg_w_param_decoder_param_latch_range427w428w(0) AND wire_w_param_decoder_param_latch_range429w(0);
	wire_w_lg_idle477w(0) <= idle AND wire_w_lg_read_param476w(0);
	wire_w_lg_read_address181w(0) <= read_address AND wire_dffe4a_w_q_range178w(0);
	wire_w_lg_read_address232w(0) <= read_address AND wire_dffe4a_w_q_range230w(0);
	wire_w_lg_read_address237w(0) <= read_address AND wire_dffe4a_w_q_range235w(0);
	wire_w_lg_read_address242w(0) <= read_address AND wire_dffe4a_w_q_range240w(0);
	wire_w_lg_read_address247w(0) <= read_address AND wire_dffe4a_w_q_range245w(0);
	wire_w_lg_read_address252w(0) <= read_address AND wire_dffe4a_w_q_range250w(0);
	wire_w_lg_read_address257w(0) <= read_address AND wire_dffe4a_w_q_range255w(0);
	wire_w_lg_read_address262w(0) <= read_address AND wire_dffe4a_w_q_range260w(0);
	wire_w_lg_read_address267w(0) <= read_address AND wire_dffe4a_w_q_range265w(0);
	wire_w_lg_read_address272w(0) <= read_address AND wire_dffe4a_w_q_range270w(0);
	wire_w_lg_read_address277w(0) <= read_address AND wire_dffe4a_w_q_range275w(0);
	wire_w_lg_read_address187w(0) <= read_address AND wire_dffe4a_w_q_range185w(0);
	wire_w_lg_read_address282w(0) <= read_address AND wire_dffe4a_w_q_range280w(0);
	wire_w_lg_read_address287w(0) <= read_address AND wire_dffe4a_w_q_range285w(0);
	wire_w_lg_read_address292w(0) <= read_address AND wire_dffe4a_w_q_range290w(0);
	wire_w_lg_read_address297w(0) <= read_address AND wire_dffe4a_w_q_range295w(0);
	wire_w_lg_read_address192w(0) <= read_address AND wire_dffe4a_w_q_range190w(0);
	wire_w_lg_read_address197w(0) <= read_address AND wire_dffe4a_w_q_range195w(0);
	wire_w_lg_read_address202w(0) <= read_address AND wire_dffe4a_w_q_range200w(0);
	wire_w_lg_read_address207w(0) <= read_address AND wire_dffe4a_w_q_range205w(0);
	wire_w_lg_read_address212w(0) <= read_address AND wire_dffe4a_w_q_range210w(0);
	wire_w_lg_read_address217w(0) <= read_address AND wire_dffe4a_w_q_range215w(0);
	wire_w_lg_read_address222w(0) <= read_address AND wire_dffe4a_w_q_range220w(0);
	wire_w_lg_read_address227w(0) <= read_address AND wire_dffe4a_w_q_range225w(0);
	wire_w_lg_read_data491w(0) <= read_data AND wire_w_lg_width_counter_param_width_match490w(0);
	wire_w_lg_read_init_counter487w(0) <= read_init_counter AND wire_w_lg_bit_counter_param_start_match485w(0);
	wire_w_lg_read_post497w(0) <= read_post AND wire_w_lg_width_counter_all_done489w(0);
	wire_w_lg_read_pre_data486w(0) <= read_pre_data AND wire_w_lg_bit_counter_param_start_match485w(0);
	wire_w_lg_rublock_regout_reg529w(0) <= rublock_regout_reg AND wire_w_lg_select_shift_nloop528w(0);
	wire_w_lg_shift_reg_load_enable77w(0) <= shift_reg_load_enable AND wire_w_data_in_range76w(0);
	wire_w_lg_shift_reg_load_enable117w(0) <= shift_reg_load_enable AND wire_w_data_in_range116w(0);
	wire_w_lg_shift_reg_load_enable121w(0) <= shift_reg_load_enable AND wire_w_data_in_range120w(0);
	wire_w_lg_shift_reg_load_enable125w(0) <= shift_reg_load_enable AND wire_w_data_in_range124w(0);
	wire_w_lg_shift_reg_load_enable129w(0) <= shift_reg_load_enable AND wire_w_data_in_range128w(0);
	wire_w_lg_shift_reg_load_enable133w(0) <= shift_reg_load_enable AND wire_w_data_in_range132w(0);
	wire_w_lg_shift_reg_load_enable137w(0) <= shift_reg_load_enable AND wire_w_data_in_range136w(0);
	wire_w_lg_shift_reg_load_enable141w(0) <= shift_reg_load_enable AND wire_w_data_in_range140w(0);
	wire_w_lg_shift_reg_load_enable145w(0) <= shift_reg_load_enable AND wire_w_data_in_range144w(0);
	wire_w_lg_shift_reg_load_enable149w(0) <= shift_reg_load_enable AND wire_w_data_in_range148w(0);
	wire_w_lg_shift_reg_load_enable153w(0) <= shift_reg_load_enable AND wire_w_data_in_range152w(0);
	wire_w_lg_shift_reg_load_enable81w(0) <= shift_reg_load_enable AND wire_w_data_in_range80w(0);
	wire_w_lg_shift_reg_load_enable157w(0) <= shift_reg_load_enable AND wire_w_data_in_range156w(0);
	wire_w_lg_shift_reg_load_enable161w(0) <= shift_reg_load_enable AND wire_w_data_in_range160w(0);
	wire_w_lg_shift_reg_load_enable165w(0) <= shift_reg_load_enable AND wire_w_data_in_range164w(0);
	wire_w_lg_shift_reg_load_enable73w(0) <= shift_reg_load_enable AND wire_w_data_in_range72w(0);
	wire_w_lg_shift_reg_load_enable85w(0) <= shift_reg_load_enable AND wire_w_data_in_range84w(0);
	wire_w_lg_shift_reg_load_enable89w(0) <= shift_reg_load_enable AND wire_w_data_in_range88w(0);
	wire_w_lg_shift_reg_load_enable93w(0) <= shift_reg_load_enable AND wire_w_data_in_range92w(0);
	wire_w_lg_shift_reg_load_enable97w(0) <= shift_reg_load_enable AND wire_w_data_in_range96w(0);
	wire_w_lg_shift_reg_load_enable101w(0) <= shift_reg_load_enable AND wire_w_data_in_range100w(0);
	wire_w_lg_shift_reg_load_enable105w(0) <= shift_reg_load_enable AND wire_w_data_in_range104w(0);
	wire_w_lg_shift_reg_load_enable109w(0) <= shift_reg_load_enable AND wire_w_data_in_range108w(0);
	wire_w_lg_shift_reg_load_enable113w(0) <= shift_reg_load_enable AND wire_w_data_in_range112w(0);
	wire_w_lg_write_data506w(0) <= write_data AND wire_w_lg_width_counter_param_width_match490w(0);
	wire_w_lg_write_init_counter503w(0) <= write_init_counter AND wire_w_lg_bit_counter_param_start_match485w(0);
	wire_w_lg_write_post_data512w(0) <= write_post_data AND wire_w_lg_bit_counter_all_done505w(0);
	wire_w_lg_write_pre_data502w(0) <= write_pre_data AND wire_w_lg_bit_counter_param_start_match485w(0);
	wire_w_lg_w_param_range173w174w(0) <= wire_w_param_range173w(0) AND wire_w_lg_w_param_range171w172w(0);
	wire_w_lg_w_param_decoder_param_latch_range427w445w(0) <= wire_w_param_decoder_param_latch_range427w(0) AND wire_w_lg_w_param_decoder_param_latch_range429w430w(0);
	wire_w_lg_w_param_decoder_param_latch_range427w440w(0) <= wire_w_param_decoder_param_latch_range427w(0) AND wire_w_param_decoder_param_latch_range429w(0);
	wire_w_lg_bit_counter_all_done505w(0) <= NOT bit_counter_all_done;
	wire_w_lg_bit_counter_param_start_match485w(0) <= NOT bit_counter_param_start_match;
	wire_w_lg_idle460w(0) <= NOT idle;
	wire_w_lg_read_address179w(0) <= NOT read_address;
	wire_w_lg_read_data456w(0) <= NOT read_data;
	wire_w_lg_read_init459w(0) <= NOT read_init;
	wire_w_lg_read_init_counter458w(0) <= NOT read_init_counter;
	wire_w_lg_read_param476w(0) <= NOT read_param;
	wire_w_lg_read_post455w(0) <= NOT read_post;
	wire_w_lg_read_pre_data457w(0) <= NOT read_pre_data;
	wire_w_lg_select_shift_nloop528w(0) <= NOT select_shift_nloop;
	wire_w_lg_shift_reg_load_enable70w(0) <= NOT shift_reg_load_enable;
	wire_w_lg_w8w168w(0) <= NOT w8w;
	wire_w_lg_width_counter_all_done489w(0) <= NOT width_counter_all_done;
	wire_w_lg_width_counter_param_width_match490w(0) <= NOT width_counter_param_width_match;
	wire_w_lg_write_data451w(0) <= NOT write_data;
	wire_w_lg_write_init454w(0) <= NOT write_init;
	wire_w_lg_write_init_counter453w(0) <= NOT write_init_counter;
	wire_w_lg_write_load449w(0) <= NOT write_load;
	wire_w_lg_write_param475w(0) <= NOT write_param;
	wire_w_lg_write_post_data450w(0) <= NOT write_post_data;
	wire_w_lg_write_pre_data452w(0) <= NOT write_pre_data;
	wire_w_lg_write_wait448w(0) <= NOT write_wait;
	wire_w_lg_w_param_range171w172w(0) <= NOT wire_w_param_range171w(0);
	wire_w_lg_w_param_decoder_param_latch_range427w428w(0) <= NOT wire_w_param_decoder_param_latch_range427w(0);
	wire_w_lg_w_param_decoder_param_latch_range429w430w(0) <= NOT wire_w_param_decoder_param_latch_range429w(0);
	wire_w_lg_w_param_decoder_param_latch_range432w433w(0) <= NOT wire_w_param_decoder_param_latch_range432w(0);
	wire_w_lg_w_lg_w_lg_idle477w478w479w(0) <= wire_w_lg_w_lg_idle477w478w(0) OR write_wait;
	wire_w_lg_w_lg_read_address181w182w(0) <= wire_w_lg_read_address181w(0) OR wire_w_lg_w_lg_read_address179w180w(0);
	wire_w_lg_w_lg_read_address232w233w(0) <= wire_w_lg_read_address232w(0) OR wire_w_lg_w_lg_read_address179w231w(0);
	wire_w_lg_w_lg_read_address237w238w(0) <= wire_w_lg_read_address237w(0) OR wire_w_lg_w_lg_read_address179w236w(0);
	wire_w_lg_w_lg_read_address242w243w(0) <= wire_w_lg_read_address242w(0) OR wire_w_lg_w_lg_read_address179w241w(0);
	wire_w_lg_w_lg_read_address247w248w(0) <= wire_w_lg_read_address247w(0) OR wire_w_lg_w_lg_read_address179w246w(0);
	wire_w_lg_w_lg_read_address252w253w(0) <= wire_w_lg_read_address252w(0) OR wire_w_lg_w_lg_read_address179w251w(0);
	wire_w_lg_w_lg_read_address257w258w(0) <= wire_w_lg_read_address257w(0) OR wire_w_lg_w_lg_read_address179w256w(0);
	wire_w_lg_w_lg_read_address262w263w(0) <= wire_w_lg_read_address262w(0) OR wire_w_lg_w_lg_read_address179w261w(0);
	wire_w_lg_w_lg_read_address267w268w(0) <= wire_w_lg_read_address267w(0) OR wire_w_lg_w_lg_read_address179w266w(0);
	wire_w_lg_w_lg_read_address272w273w(0) <= wire_w_lg_read_address272w(0) OR wire_w_lg_w_lg_read_address179w271w(0);
	wire_w_lg_w_lg_read_address277w278w(0) <= wire_w_lg_read_address277w(0) OR wire_w_lg_w_lg_read_address179w276w(0);
	wire_w_lg_w_lg_read_address187w188w(0) <= wire_w_lg_read_address187w(0) OR wire_w_lg_w_lg_read_address179w186w(0);
	wire_w_lg_w_lg_read_address282w283w(0) <= wire_w_lg_read_address282w(0) OR wire_w_lg_w_lg_read_address179w281w(0);
	wire_w_lg_w_lg_read_address287w288w(0) <= wire_w_lg_read_address287w(0) OR wire_w_lg_w_lg_read_address179w286w(0);
	wire_w_lg_w_lg_read_address292w293w(0) <= wire_w_lg_read_address292w(0) OR wire_w_lg_w_lg_read_address179w291w(0);
	wire_w_lg_w_lg_read_address297w298w(0) <= wire_w_lg_read_address297w(0) OR wire_w_lg_w_lg_read_address179w296w(0);
	wire_w_lg_w_lg_read_address192w193w(0) <= wire_w_lg_read_address192w(0) OR wire_w_lg_w_lg_read_address179w191w(0);
	wire_w_lg_w_lg_read_address197w198w(0) <= wire_w_lg_read_address197w(0) OR wire_w_lg_w_lg_read_address179w196w(0);
	wire_w_lg_w_lg_read_address202w203w(0) <= wire_w_lg_read_address202w(0) OR wire_w_lg_w_lg_read_address179w201w(0);
	wire_w_lg_w_lg_read_address207w208w(0) <= wire_w_lg_read_address207w(0) OR wire_w_lg_w_lg_read_address179w206w(0);
	wire_w_lg_w_lg_read_address212w213w(0) <= wire_w_lg_read_address212w(0) OR wire_w_lg_w_lg_read_address179w211w(0);
	wire_w_lg_w_lg_read_address217w218w(0) <= wire_w_lg_read_address217w(0) OR wire_w_lg_w_lg_read_address179w216w(0);
	wire_w_lg_w_lg_read_address222w223w(0) <= wire_w_lg_read_address222w(0) OR wire_w_lg_w_lg_read_address179w221w(0);
	wire_w_lg_w_lg_read_address227w228w(0) <= wire_w_lg_read_address227w(0) OR wire_w_lg_w_lg_read_address179w226w(0);
	wire_w_lg_w_lg_shift_reg_load_enable67w68w(0) <= wire_w_lg_shift_reg_load_enable67w(0) OR shift_reg_clear;
	wire_w_lg_shift_reg_load_enable67w(0) <= shift_reg_load_enable OR shift_reg_shift_enable;
	bit_counter_all_done <= (((((wire_cntr2_q(0) AND wire_cntr2_q(1)) AND (NOT wire_cntr2_q(2))) AND wire_cntr2_q(3)) AND (NOT wire_cntr2_q(4))) AND wire_cntr2_q(5));
	bit_counter_clear <= (read_init OR write_init);
	bit_counter_enable <= (((((((((read_init OR write_init) OR read_init_counter) OR write_init_counter) OR read_pre_data) OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data);
	bit_counter_param_start <= start_bit_decoder_out;
	bit_counter_param_start_match <= ((((((NOT w22w(0)) AND (NOT w22w(1))) AND (NOT w22w(2))) AND (NOT w22w(3))) AND (NOT w22w(4))) AND (NOT w22w(5)));
	busy <= wire_w_lg_idle460w(0);
	data_out <= ( wire_w_lg_w_lg_read_address297w298w & wire_w_lg_w_lg_read_address292w293w & wire_w_lg_w_lg_read_address287w288w & wire_w_lg_w_lg_read_address282w283w & wire_w_lg_w_lg_read_address277w278w & wire_w_lg_w_lg_read_address272w273w & wire_w_lg_w_lg_read_address267w268w & wire_w_lg_w_lg_read_address262w263w & wire_w_lg_w_lg_read_address257w258w & wire_w_lg_w_lg_read_address252w253w & wire_w_lg_w_lg_read_address247w248w & wire_w_lg_w_lg_read_address242w243w & wire_w_lg_w_lg_read_address237w238w & wire_w_lg_w_lg_read_address232w233w & wire_w_lg_w_lg_read_address227w228w & wire_w_lg_w_lg_read_address222w223w & wire_w_lg_w_lg_read_address217w218w & wire_w_lg_w_lg_read_address212w213w & wire_w_lg_w_lg_read_address207w208w & wire_w_lg_w_lg_read_address202w203w & wire_w_lg_w_lg_read_address197w198w & wire_w_lg_w_lg_read_address192w193w & wire_w_lg_w_lg_read_address187w188w & wire_w_lg_w_lg_read_address181w182w);
	idle <= idle_state;
	param_decoder_param_latch <= dffe6a;
	param_decoder_select <= ( wire_w446w & wire_w_lg_w431w443w & wire_w441w & wire_w_lg_w437w438w & wire_w_lg_w431w434w);
	power_up <= ((((((((((((wire_w_lg_idle460w(0) AND wire_w_lg_read_init459w(0)) AND wire_w_lg_read_init_counter458w(0)) AND wire_w_lg_read_pre_data457w(0)) AND wire_w_lg_read_data456w(0)) AND wire_w_lg_read_post455w(0)) AND wire_w_lg_write_init454w(0)) AND wire_w_lg_write_init_counter453w(0)) AND wire_w_lg_write_pre_data452w(0)) AND wire_w_lg_write_data451w(0)) AND wire_w_lg_write_post_data450w(0)) AND wire_w_lg_write_load449w(0)) AND wire_w_lg_write_wait448w(0));
	read_address <= read_address_state;
	read_data <= read_data_state;
	read_init <= read_init_state;
	read_init_counter <= read_init_counter_state;
	read_post <= read_post_state;
	read_pre_data <= read_pre_data_state;
	rublock_captnupdt <= wire_w_lg_write_load449w(0);
	rublock_clock <= (NOT (clock OR idle_write_wait));
	rublock_reconfig <= rublock_reconfig_st;
	rublock_reconfig_st <= (idle AND reconfig);
	rublock_regin <= (wire_w_lg_rublock_regout_reg529w(0) OR (shift_reg_serial_out AND select_shift_nloop));
	rublock_regout <= wire_sd1_regout;
	rublock_regout_reg <= dffe5;
	rublock_shiftnld <= (((((read_pre_data OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data);
	select_shift_nloop <= (wire_w_lg_read_data491w(0) OR wire_w_lg_write_data506w(0));
	shift_reg_clear <= read_init;
	shift_reg_load_enable <= (idle AND write_param);
	shift_reg_serial_in <= (rublock_regout_reg AND select_shift_nloop);
	shift_reg_serial_out <= dffe4a(0);
	shift_reg_shift_enable <= (((read_data OR write_data) OR read_post) OR write_post_data);
	start_bit_decoder_out <= ((((( "0" & "0" & "0" & "0" & "0" & "0") OR ( "0" & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1))) OR ( "0" & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & "0")) OR ( "0" & "0" & "0" & start_bit_decoder_param_select(3) & start_bit_decoder_param_select(3) & "0")) OR ( "0" & "0" & "0" & start_bit_decoder_param_select(4) & "0" & start_bit_decoder_param_select(4)));
	start_bit_decoder_param_select <= param_decoder_select;
	w22w <= (wire_cntr2_q XOR bit_counter_param_start);
	w51w <= (wire_cntr3_q XOR width_counter_param_width);
	w8w <= wire_w_lg_idle460w(0);
	width_counter_all_done <= ((((wire_cntr3_q(0) AND wire_cntr3_q(1)) AND wire_cntr3_q(2)) AND (NOT wire_cntr3_q(3))) AND wire_cntr3_q(4));
	width_counter_clear <= (read_init OR write_init);
	width_counter_enable <= ((read_data OR write_data) OR read_post);
	width_counter_param_width <= width_decoder_out;
	width_counter_param_width_match <= (((((NOT w51w(0)) AND (NOT w51w(1))) AND (NOT w51w(2))) AND (NOT w51w(3))) AND (NOT w51w(4)));
	width_decoder_out <= ((((( "0" & "0" & width_decoder_param_select(0) & "0" & width_decoder_param_select(0)) OR ( "0" & width_decoder_param_select(1) & width_decoder_param_select(1) & "0" & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(2))) OR ( width_decoder_param_select(3) & width_decoder_param_select(3) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(4)));
	width_decoder_param_select <= param_decoder_select;
	write_data <= write_data_state;
	write_init <= write_init_state;
	write_init_counter <= write_init_counter_state;
	write_load <= write_load_state;
	write_post_data <= write_post_data_state;
	write_pre_data <= write_pre_data_state;
	write_wait <= write_wait_state;
	wire_w_data_in_range76w(0) <= data_in(0);
	wire_w_data_in_range116w(0) <= data_in(10);
	wire_w_data_in_range120w(0) <= data_in(11);
	wire_w_data_in_range124w(0) <= data_in(12);
	wire_w_data_in_range128w(0) <= data_in(13);
	wire_w_data_in_range132w(0) <= data_in(14);
	wire_w_data_in_range136w(0) <= data_in(15);
	wire_w_data_in_range140w(0) <= data_in(16);
	wire_w_data_in_range144w(0) <= data_in(17);
	wire_w_data_in_range148w(0) <= data_in(18);
	wire_w_data_in_range152w(0) <= data_in(19);
	wire_w_data_in_range80w(0) <= data_in(1);
	wire_w_data_in_range156w(0) <= data_in(20);
	wire_w_data_in_range160w(0) <= data_in(21);
	wire_w_data_in_range164w(0) <= data_in(22);
	wire_w_data_in_range72w(0) <= data_in(23);
	wire_w_data_in_range84w(0) <= data_in(2);
	wire_w_data_in_range88w(0) <= data_in(3);
	wire_w_data_in_range92w(0) <= data_in(4);
	wire_w_data_in_range96w(0) <= data_in(5);
	wire_w_data_in_range100w(0) <= data_in(6);
	wire_w_data_in_range104w(0) <= data_in(7);
	wire_w_data_in_range108w(0) <= data_in(8);
	wire_w_data_in_range112w(0) <= data_in(9);
	wire_w_param_range171w(0) <= param(1);
	wire_w_param_range173w(0) <= param(2);
	wire_w_param_decoder_param_latch_range427w(0) <= param_decoder_param_latch(0);
	wire_w_param_decoder_param_latch_range429w(0) <= param_decoder_param_latch(1);
	wire_w_param_decoder_param_latch_range432w(0) <= param_decoder_param_latch(2);
	check_busy_dffe <= (OTHERS => '0');
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(0) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(0) <= '0';
				ELSE dffe4a(0) <= (wire_w_lg_shift_reg_load_enable77w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w75w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(1) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(1) <= '0';
				ELSE dffe4a(1) <= (wire_w_lg_shift_reg_load_enable81w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w79w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(2) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(2) <= '0';
				ELSE dffe4a(2) <= (wire_w_lg_shift_reg_load_enable85w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w83w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(3) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(3) <= '0';
				ELSE dffe4a(3) <= (wire_w_lg_shift_reg_load_enable89w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w87w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(4) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(4) <= '0';
				ELSE dffe4a(4) <= (wire_w_lg_shift_reg_load_enable93w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w91w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(5) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(5) <= '0';
				ELSE dffe4a(5) <= (wire_w_lg_shift_reg_load_enable97w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w95w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(6) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(6) <= '0';
				ELSE dffe4a(6) <= (wire_w_lg_shift_reg_load_enable101w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w99w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(7) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(7) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(7) <= '0';
				ELSE dffe4a(7) <= (wire_w_lg_shift_reg_load_enable105w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w103w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(8) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(8) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(8) <= '0';
				ELSE dffe4a(8) <= (wire_w_lg_shift_reg_load_enable109w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w107w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(9) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(9) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(9) <= '0';
				ELSE dffe4a(9) <= (wire_w_lg_shift_reg_load_enable113w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w111w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(10) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(10) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(10) <= '0';
				ELSE dffe4a(10) <= (wire_w_lg_shift_reg_load_enable117w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w115w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(11) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(11) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(11) <= '0';
				ELSE dffe4a(11) <= (wire_w_lg_shift_reg_load_enable121w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w119w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(12) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(12) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(12) <= '0';
				ELSE dffe4a(12) <= (wire_w_lg_shift_reg_load_enable125w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w123w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(13) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(13) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(13) <= '0';
				ELSE dffe4a(13) <= (wire_w_lg_shift_reg_load_enable129w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w127w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(14) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(14) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(14) <= '0';
				ELSE dffe4a(14) <= (wire_w_lg_shift_reg_load_enable133w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w131w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(15) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(15) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(15) <= '0';
				ELSE dffe4a(15) <= (wire_w_lg_shift_reg_load_enable137w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w135w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(16) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(16) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(16) <= '0';
				ELSE dffe4a(16) <= (wire_w_lg_shift_reg_load_enable141w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w139w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(17) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(17) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(17) <= '0';
				ELSE dffe4a(17) <= (wire_w_lg_shift_reg_load_enable145w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w143w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(18) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(18) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(18) <= '0';
				ELSE dffe4a(18) <= (wire_w_lg_shift_reg_load_enable149w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w147w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(19) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(19) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(19) <= '0';
				ELSE dffe4a(19) <= (wire_w_lg_shift_reg_load_enable153w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w151w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(20) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(20) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(20) <= '0';
				ELSE dffe4a(20) <= (wire_w_lg_shift_reg_load_enable157w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w155w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(21) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(21) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(21) <= '0';
				ELSE dffe4a(21) <= (wire_w_lg_shift_reg_load_enable161w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w159w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(22) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(22) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(22) <= '0';
				ELSE dffe4a(22) <= (wire_w_lg_shift_reg_load_enable165w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w163w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe4a(23) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ena(23) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe4a(23) <= '0';
				ELSE dffe4a(23) <= (wire_w_lg_shift_reg_load_enable73w(0) OR wire_w_lg_w_lg_shift_reg_load_enable70w71w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	loop0 : FOR i IN 0 TO 23 GENERATE
		wire_dffe4a_ena(i) <= wire_w_lg_w_lg_shift_reg_load_enable67w68w(0);
	END GENERATE loop0;
	wire_dffe4a_w_q_range178w(0) <= dffe4a(0);
	wire_dffe4a_w_q_range230w(0) <= dffe4a(10);
	wire_dffe4a_w_q_range235w(0) <= dffe4a(11);
	wire_dffe4a_w_q_range240w(0) <= dffe4a(12);
	wire_dffe4a_w_q_range245w(0) <= dffe4a(13);
	wire_dffe4a_w_q_range250w(0) <= dffe4a(14);
	wire_dffe4a_w_q_range255w(0) <= dffe4a(15);
	wire_dffe4a_w_q_range260w(0) <= dffe4a(16);
	wire_dffe4a_w_q_range265w(0) <= dffe4a(17);
	wire_dffe4a_w_q_range270w(0) <= dffe4a(18);
	wire_dffe4a_w_q_range275w(0) <= dffe4a(19);
	wire_dffe4a_w_q_range185w(0) <= dffe4a(1);
	wire_dffe4a_w_q_range280w(0) <= dffe4a(20);
	wire_dffe4a_w_q_range285w(0) <= dffe4a(21);
	wire_dffe4a_w_q_range290w(0) <= dffe4a(22);
	wire_dffe4a_w_q_range295w(0) <= dffe4a(23);
	wire_dffe4a_w_q_range190w(0) <= dffe4a(2);
	wire_dffe4a_w_q_range195w(0) <= dffe4a(3);
	wire_dffe4a_w_q_range200w(0) <= dffe4a(4);
	wire_dffe4a_w_q_range205w(0) <= dffe4a(5);
	wire_dffe4a_w_q_range210w(0) <= dffe4a(6);
	wire_dffe4a_w_q_range215w(0) <= dffe4a(7);
	wire_dffe4a_w_q_range220w(0) <= dffe4a(8);
	wire_dffe4a_w_q_range225w(0) <= dffe4a(9);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe5 <= rublock_regout;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe6a(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe6a_ena(0) = '1') THEN dffe6a(0) <= param(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe6a(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe6a_ena(1) = '1') THEN dffe6a(1) <= param(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe6a(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe6a_ena(2) = '1') THEN dffe6a(2) <= param(2);
			END IF;
		END IF;
	END PROCESS;
	loop1 : FOR i IN 0 TO 2 GENERATE
		wire_dffe6a_ena(i) <= (idle AND (write_param OR read_param));
	END GENERATE loop1;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN idle_state <= '1';
		ELSIF (clock = '1' AND clock'event) THEN idle_state <= (((wire_w_lg_w_lg_w_lg_idle477w478w479w(0) OR (read_data AND width_counter_all_done)) OR (read_post AND width_counter_all_done)) OR power_up);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN idle_write_wait <= '0';
		ELSIF (clock = '1' AND clock'event) THEN idle_write_wait <= ((((wire_w_lg_w_lg_w_lg_idle477w478w479w(0) OR (read_data AND width_counter_all_done)) OR (read_post AND width_counter_all_done)) OR power_up) AND write_load);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_address_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_read_address_state_ena = '1') THEN read_address_state <= (((read_param OR write_param) AND (wire_w_lg_w_param_range173w174w(0) AND (NOT param(0)))) AND wire_w_lg_w8w168w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_read_address_state_ena <= (read_param OR write_param);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_data_state <= (((read_init_counter AND bit_counter_param_start_match) OR (read_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_read_data491w(0) AND wire_w_lg_width_counter_all_done489w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_init_counter_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_init_counter_state <= read_init;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_init_state <= (idle AND read_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_post_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_post_state <= (((read_data AND width_counter_param_width_match) AND wire_w_lg_width_counter_all_done489w(0)) OR wire_w_lg_read_post497w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_pre_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_pre_data_state <= (wire_w_lg_read_init_counter487w(0) OR wire_w_lg_read_pre_data486w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_data_state <= (((write_init_counter AND bit_counter_param_start_match) OR (write_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_write_data506w(0) AND wire_w_lg_bit_counter_all_done505w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_init_counter_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_init_counter_state <= write_init;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_init_state <= (idle AND write_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_load_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_load_state <= ((write_data AND bit_counter_all_done) OR (write_post_data AND bit_counter_all_done));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_post_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_post_data_state <= (((write_data AND width_counter_param_width_match) AND wire_w_lg_bit_counter_all_done505w(0)) OR wire_w_lg_write_post_data512w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_pre_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_pre_data_state <= (wire_w_lg_write_init_counter503w(0) OR wire_w_lg_write_pre_data502w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_wait_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_wait_state <= write_load;
		END IF;
	END PROCESS;
	cntr2 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		aclr => reset,
		clock => clock,
		cnt_en => bit_counter_enable,
		q => wire_cntr2_q,
		sclr => bit_counter_clear
	  );
	cntr3 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		aclr => reset,
		clock => clock,
		cnt_en => width_counter_enable,
		q => wire_cntr3_q,
		sclr => width_counter_clear
	  );
	sd1 :  arriaii_rublock
	  PORT MAP ( 
		captnupdt => rublock_captnupdt,
		clk => rublock_clock,
		rconfig => rublock_reconfig,
		regin => rublock_regin,
		regout => wire_sd1_regout,
		rsttimer => reset_timer,
		shiftnld => rublock_shiftnld
	  );

 END RTL; --remote_update_rmtupdt_6co
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY remote_update IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data_in		: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		param		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		read_param		: IN STD_LOGIC ;
		reconfig		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		reset_timer		: IN STD_LOGIC ;
		write_param		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_out		: OUT STD_LOGIC_VECTOR (23 DOWNTO 0)
	);
END remote_update;


ARCHITECTURE RTL OF remote_update IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "altremote_update";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "check_app_pof=false;config_device_addr_width=24;intended_device_family=Arria II GX;in_data_width=24;operation_mode=REMOTE;out_data_width=24;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (23 DOWNTO 0);



	COMPONENT remote_update_rmtupdt_6co
	PORT (
			clock	: IN STD_LOGIC ;
			data_in	: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
			read_param	: IN STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			data_out	: OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
			param	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig	: IN STD_LOGIC ;
			reset	: IN STD_LOGIC ;
			reset_timer	: IN STD_LOGIC ;
			write_param	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	busy    <= sub_wire0;
	data_out    <= sub_wire1(23 DOWNTO 0);

	remote_update_rmtupdt_6co_component : remote_update_rmtupdt_6co
	PORT MAP (
		clock => clock,
		data_in => data_in,
		read_param => read_param,
		param => param,
		reconfig => reconfig,
		reset => reset,
		reset_timer => reset_timer,
		write_param => write_param,
		busy => sub_wire0,
		data_out => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: PRIVATE: SIM_INIT_PAGE_SELECT_COMBO STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT0_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT1_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT2_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT3_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT4_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_WATCHDOG_VALUE_EDIT STRING "1"
-- Retrieval info: PRIVATE: SUPPORT_WRITE_CHECK STRING "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WATCHDOG_ENABLE_CHECK STRING "0"
-- Retrieval info: CONSTANT: CHECK_APP_POF STRING "false"
-- Retrieval info: CONSTANT: CONFIG_DEVICE_ADDR_WIDTH NUMERIC "24"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: CONSTANT: IN_DATA_WIDTH NUMERIC "24"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "REMOTE"
-- Retrieval info: CONSTANT: OUT_DATA_WIDTH NUMERIC "24"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data_in 0 0 24 0 INPUT NODEFVAL "data_in[23..0]"
-- Retrieval info: USED_PORT: data_out 0 0 24 0 OUTPUT NODEFVAL "data_out[23..0]"
-- Retrieval info: USED_PORT: param 0 0 3 0 INPUT NODEFVAL "param[2..0]"
-- Retrieval info: USED_PORT: read_param 0 0 0 0 INPUT NODEFVAL "read_param"
-- Retrieval info: USED_PORT: reconfig 0 0 0 0 INPUT NODEFVAL "reconfig"
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: USED_PORT: reset_timer 0 0 0 0 INPUT NODEFVAL "reset_timer"
-- Retrieval info: USED_PORT: write_param 0 0 0 0 INPUT NODEFVAL "write_param"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data_in 0 0 24 0 data_in 0 0 24 0
-- Retrieval info: CONNECT: @param 0 0 3 0 param 0 0 3 0
-- Retrieval info: CONNECT: @read_param 0 0 0 0 read_param 0 0 0 0
-- Retrieval info: CONNECT: @reconfig 0 0 0 0 reconfig 0 0 0 0
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: CONNECT: @reset_timer 0 0 0 0 reset_timer 0 0 0 0
-- Retrieval info: CONNECT: @write_param 0 0 0 0 write_param 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: data_out 0 0 24 0 @data_out 0 0 24 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update_inst.vhd FALSE
-- Retrieval info: LIB_FILE: arriaii
-- Retrieval info: LIB_FILE: lpm
