-- megafunction wizard: %ALTASMI_PARALLEL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTASMI_PARALLEL 

-- ============================================================
-- File Name: altasmi.vhd
-- Megafunction Name(s):
-- 			ALTASMI_PARALLEL
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altasmi_parallel CBX_AUTO_BLACKBOX="ALL" DATA_WIDTH="STANDARD" DEVICE_FAMILY="Arria II GX" EPCS_TYPE="EPCS128" PAGE_SIZE=256 PORT_BULK_ERASE="PORT_UNUSED" PORT_DIE_ERASE="PORT_UNUSED" PORT_EN4B_ADDR="PORT_UNUSED" PORT_EX4B_ADDR="PORT_UNUSED" PORT_FAST_READ="PORT_USED" PORT_ILLEGAL_ERASE="PORT_USED" PORT_ILLEGAL_WRITE="PORT_USED" PORT_RDID_OUT="PORT_USED" PORT_READ_ADDRESS="PORT_USED" PORT_READ_DUMMYCLK="PORT_UNUSED" PORT_READ_RDID="PORT_USED" PORT_READ_SID="PORT_UNUSED" PORT_READ_STATUS="PORT_USED" PORT_SECTOR_ERASE="PORT_USED" PORT_SECTOR_PROTECT="PORT_UNUSED" PORT_SHIFT_BYTES="PORT_USED" PORT_WREN="PORT_UNUSED" PORT_WRITE="PORT_USED" USE_ASMIBLOCK="OFF" USE_EAB="ON" WRITE_DUMMY_CLK=0 addr asmi_dataoe asmi_dataout asmi_dclk asmi_scein asmi_sdoin busy clkin data_valid datain dataout fast_read illegal_erase illegal_write rden rdid_out read_address read_rdid read_status reset sector_erase shift_bytes status_out write INTENDED_DEVICE_FAMILY="Arria II GX" ALTERA_INTERNAL_OPTIONS=SUPPRESS_DA_RULE_INTERNAL=C106
--VERSION_BEGIN 13.1 cbx_a_gray2bin 2013:10:17:04:07:49:SJ cbx_a_graycounter 2013:10:17:04:07:49:SJ cbx_altasmi_parallel 2013:10:17:04:07:49:SJ cbx_altdpram 2013:10:17:04:07:49:SJ cbx_altsyncram 2013:10:17:04:07:49:SJ cbx_arriav 2013:10:17:04:07:49:SJ cbx_cyclone 2013:10:17:04:07:49:SJ cbx_cycloneii 2013:10:17:04:07:49:SJ cbx_fifo_common 2013:10:17:04:07:49:SJ cbx_lpm_add_sub 2013:10:17:04:07:49:SJ cbx_lpm_compare 2013:10:17:04:07:49:SJ cbx_lpm_counter 2013:10:17:04:07:49:SJ cbx_lpm_decode 2013:10:17:04:07:49:SJ cbx_lpm_mux 2013:10:17:04:07:49:SJ cbx_mgl 2013:10:17:04:34:36:SJ cbx_nightfury 2013:10:17:04:07:49:SJ cbx_scfifo 2013:10:17:04:07:49:SJ cbx_stratix 2013:10:17:04:07:49:SJ cbx_stratixii 2013:10:17:04:07:49:SJ cbx_stratixiii 2013:10:17:04:07:49:SJ cbx_stratixv 2013:10:17:04:07:49:SJ cbx_util_mgl 2013:10:17:04:07:49:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = a_graycounter 4 lpm_compare 2 lpm_counter 3 lut 29 mux21 2 reg 153 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altasmi_altasmi_parallel_pu03 IS 
	 PORT 
	 ( 
		 addr	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 asmi_dataoe	:	OUT  STD_LOGIC;
		 asmi_dataout	:	IN  STD_LOGIC := '0';
		 asmi_dclk	:	OUT  STD_LOGIC;
		 asmi_scein	:	OUT  STD_LOGIC;
		 asmi_sdoin	:	OUT  STD_LOGIC;
		 busy	:	OUT  STD_LOGIC;
		 clkin	:	IN  STD_LOGIC;
		 data_valid	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 fast_read	:	IN  STD_LOGIC := '0';
		 illegal_erase	:	OUT  STD_LOGIC;
		 illegal_write	:	OUT  STD_LOGIC;
		 rden	:	IN  STD_LOGIC;
		 rdid_out	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 read_address	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 read_rdid	:	IN  STD_LOGIC := '0';
		 read_status	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC := '0';
		 sector_erase	:	IN  STD_LOGIC := '0';
		 shift_bytes	:	IN  STD_LOGIC := '0';
		 status_out	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 write	:	IN  STD_LOGIC := '0'
	 ); 
 END altasmi_altasmi_parallel_pu03;

 ARCHITECTURE RTL OF altasmi_altasmi_parallel_pu03 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "SUPPRESS_DA_RULE_INTERNAL=C106";

	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range175w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range178w179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_addbyte_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_end_operation107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range119w120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range117w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_in_operation47w48w49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_end1_cyc_reg_in_wire50w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w347w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range109w112w344w345w346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range109w112w349w350w351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range109w110w111w358w359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w114w435w436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w112w344w345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w112w369w370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w112w349w350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w110w111w358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range109w114w435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range109w112w344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range109w112w369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range109w112w349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range109w112w171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range109w112w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range108w113w139w140w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range108w113w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range109w110w111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range109w114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range109w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range108w113w139w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range108w113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range109w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w103w104w105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w_q_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_q_range109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_lg_w_q_range638w639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_lg_w_q_range636w637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w631w632w633w634w635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_wrstage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_q_range636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_q_range638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 add_msb_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_add_msb_reg_ena	:	STD_LOGIC;
	 SIGNAL	 add_rollover_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 addr_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range408w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_asmi_opcode_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 asmi_opcode_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_asmi_opcode_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_asmi_opcode_reg_w_q_range185w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 buf_empty_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 busy_delay_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 busy_det_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rdid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rstat_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_write_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cnt_bfend_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 do_wrmemadd_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dvalid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dvalid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_dvalid_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 dvalid_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_hdlyreg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_pgwrop_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_pgwrop_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_rbyte_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_rbyte_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_end_rbyte_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 end_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 fast_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_fast_read_reg_ena	:	STD_LOGIC;
	 SIGNAL	 ill_erase_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ill_write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 illegal_erase_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 illegal_write_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 illegal_write_prot_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_cnt_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 maxcnt_shift_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 maxcnt_shift_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ncs_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_ncs_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_ncs_reg_w_lg_q395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_pgwrbuf_dataout_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 pgwrbuf_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_pgwrbuf_dataout_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_pgwrbuf_dataout_w_q_range579w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 power_up_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rdid_out_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_add_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 read_add_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_add_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL	 read_bufdly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_data_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_read_dout_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_dout_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_dout_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 read_rdid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_rdid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 read_status_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_status_reg_ena	:	STD_LOGIC;
	 SIGNAL	 sec_erase_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_sec_erase_reg_ena	:	STD_LOGIC;
	 SIGNAL	 shftpgwr_data_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage2_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage4_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 start_wrpoll_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_start_wrpoll_reg_ena	:	STD_LOGIC;
	 SIGNAL	 start_wrpoll_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_int_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 statreg_int	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_int_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_statreg_out_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 statreg_out	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_out_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 write_prot_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_write_prot_reg_ena	:	STD_LOGIC;
	 SIGNAL	 write_prot_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_write_reg_ena	:	STD_LOGIC;
	 SIGNAL	 write_rstat_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cmpr4_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr4_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr4_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr5_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr5_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_q	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_read_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_read_buf774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_read_cntr_q	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire498w499w500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_data	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_q	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_rden_wire498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	wire_mux211_dataout	:	STD_LOGIC;
	 SIGNAL	wire_mux212_dataout	:	STD_LOGIC;
	 SIGNAL  wire_scfifo3_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_scfifo3_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_scfifo3_rdreq	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_read_buf576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_scfifo3_wrreq	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_shift_bytes_wire574w575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_scfifo3_w_q_range582w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_scfifo3_w_q_range587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w549w550w551w552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w549w550w551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w799w800w801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w549w550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w799w800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w244w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w237w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_end_operation545w546w547w548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode201w202w203w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode201w202w203w204w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode206w207w208w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode206w207w208w209w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode240w241w242w243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode211w212w213w292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode211w212w213w214w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode252w253w254w310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode252w253w254w255w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode233w234w235w236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read374w375w376w377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write544w796w797w798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w644w791w792w802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read422w489w490w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase61w431w432w433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_end_operation545w546w547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode201w202w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode206w207w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode216w221w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode216w221w222w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode216w217w294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode216w217w218w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode240w241w242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode211w212w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode252w253w254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode233w234w235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp2_wire660w661w662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp2_wire660w661w665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp2_wire660w667w668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp2_wire660w667w670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read374w375w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read374w375w434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write544w796w797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w644w791w792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read422w489w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_erase61w431w432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire672w673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire672w675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire677w678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire677w680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_4baddr193w194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_ex4baddr188w189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_polling558w559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat129w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write224w225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write70w353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_operation545w546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_read_byte496w508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode195w284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode195w196w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode190w282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode190w191w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode226w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode226w227w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode201w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode206w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode246w306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode246w247w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode249w308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode249w250w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode229w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode229w230w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode257w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode257w258w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode260w314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode260w261w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode216w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode216w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode240w241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode211w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode252w253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode198w286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode198w199w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode233w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_reach_max_cnt626w627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage3_wire52w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_start_poll360w361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire660w661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire660w667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read374w375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write544w796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly580w581w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w631w632w633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w644w791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write79w80w423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read422w489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_rdid131w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase61w431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_operation560w561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rden_wire427w428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie407w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp2_wire672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp2_wire677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_nonvolatile340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read_byte496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy411w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_reach_max_cnt626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly583w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_opcode186w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire409w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_start_poll360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range682w695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range685w702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range687w707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range689w712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range691w717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range693w721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write70w372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w125w126w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp0_wire658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp1_wire659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp2_wire660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_buf_empty765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_busy_wire3w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clkin_wire45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_die_erase542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_fast_read373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_memadd440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_volatile232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_prot540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write_volatile239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_add_cycle90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_fast_read84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_ophdly46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_pgwr_data69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reach_max_cnt590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_rdid_wire12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_sid_wire11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_status_wire26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sec_protect_wire10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_st_busy_wire133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_start_poll128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_prot_true629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_wire20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range75w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w644w791w792w802w803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode260w314w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode260w261w262w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write79w80w423w424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_end_operation560w561w562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire427w428w429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy419w420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy411w412w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly583w584w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire458w459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode260w314w315w316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode260w261w262w263w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w631w632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_rden_wire427w428w429w430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_not_busy411w412w413w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w264w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w317w318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w264w265w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w317w318w319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w264w265w266w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w317w318w319w320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w264w265w266w267w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w317w318w319w320w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w264w265w266w267w268w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w317w318w319w320w321w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w264w265w266w267w268w269w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w270w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w323w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w270w271w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w323w324w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w270w271w272w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w323w324w325w326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w270w271w272w273w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w323w324w325w326w327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w270w271w272w273w274w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w323w324w325w326w327w328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w270w271w272w273w274w275w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w276w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w329w330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w276w277w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w276w277w278w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w168w169w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w168w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w125w126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w690w692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read422w443w444w445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read_sid164w165w166w167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bp3_wire653w654w655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read422w443w444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_sid164w165w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_stat453w454w455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_erase646w647w648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write79w122w123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_prot_wire_range666w684w686w688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp3_wire653w654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read422w457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read422w443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_sid164w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat453w454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase646w647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write79w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write79w80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly577w578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_prot_wire_range666w684w686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp3_wire653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data0out_wire461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_sid164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range703w731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range708w735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range713w739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range718w743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_add_range722w747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range705w729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range710w733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range715w737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range720w741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_check_range724w745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range595w598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range599w601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range602w604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range605w607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range608w610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range611w613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range614w616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range617w619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_prot_wire_range666w684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range682w698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range685w704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range687w709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range689w714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range691w719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mask_prot_range693w723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  add_rollover :	STD_LOGIC;
	 SIGNAL  addr_overdie :	STD_LOGIC;
	 SIGNAL  addr_overdie_pos :	STD_LOGIC;
	 SIGNAL  addr_reg_overdie :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  b4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  be_write_prot :	STD_LOGIC;
	 SIGNAL  berase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  bp0_wire :	STD_LOGIC;
	 SIGNAL  bp1_wire :	STD_LOGIC;
	 SIGNAL  bp2_wire :	STD_LOGIC;
	 SIGNAL  bp3_wire :	STD_LOGIC;
	 SIGNAL  buf_empty :	STD_LOGIC;
	 SIGNAL  busy_wire :	STD_LOGIC;
	 SIGNAL  clkin_wire :	STD_LOGIC;
	 SIGNAL  clr_addmsb_wire :	STD_LOGIC;
	 SIGNAL  clr_endrbyte_wire :	STD_LOGIC;
	 SIGNAL  clr_rdid_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire2 :	STD_LOGIC;
	 SIGNAL  clr_rstat_wire :	STD_LOGIC;
	 SIGNAL  clr_write_wire :	STD_LOGIC;
	 SIGNAL  clr_write_wire2 :	STD_LOGIC;
	 SIGNAL  cnt_bfend_wire_in :	STD_LOGIC;
	 SIGNAL  data0out_wire :	STD_LOGIC;
	 SIGNAL  data_valid_wire :	STD_LOGIC;
	 SIGNAL  dataout_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  derase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  do_4baddr :	STD_LOGIC;
	 SIGNAL  do_bulk_erase :	STD_LOGIC;
	 SIGNAL  do_die_erase :	STD_LOGIC;
	 SIGNAL  do_ex4baddr :	STD_LOGIC;
	 SIGNAL  do_fast_read :	STD_LOGIC;
	 SIGNAL  do_fread_epcq :	STD_LOGIC;
	 SIGNAL  do_freadwrv_polling :	STD_LOGIC;
	 SIGNAL  do_memadd :	STD_LOGIC;
	 SIGNAL  do_polling :	STD_LOGIC;
	 SIGNAL  do_read :	STD_LOGIC;
	 SIGNAL  do_read_nonvolatile :	STD_LOGIC;
	 SIGNAL  do_read_rdid :	STD_LOGIC;
	 SIGNAL  do_read_sid :	STD_LOGIC;
	 SIGNAL  do_read_stat :	STD_LOGIC;
	 SIGNAL  do_read_volatile :	STD_LOGIC;
	 SIGNAL  do_sec_erase :	STD_LOGIC;
	 SIGNAL  do_sec_prot :	STD_LOGIC;
	 SIGNAL  do_secprot_wren :	STD_LOGIC;
	 SIGNAL  do_sprot_polling :	STD_LOGIC;
	 SIGNAL  do_sprot_rstat :	STD_LOGIC;
	 SIGNAL  do_wait_dummyclk :	STD_LOGIC;
	 SIGNAL  do_wren :	STD_LOGIC;
	 SIGNAL  do_write :	STD_LOGIC;
	 SIGNAL  do_write_polling :	STD_LOGIC;
	 SIGNAL  do_write_rstat :	STD_LOGIC;
	 SIGNAL  do_write_volatile :	STD_LOGIC;
	 SIGNAL  do_write_volatile_rstat :	STD_LOGIC;
	 SIGNAL  do_write_volatile_wren :	STD_LOGIC;
	 SIGNAL  do_write_wren :	STD_LOGIC;
	 SIGNAL  dummy_read_buf :	STD_LOGIC;
	 SIGNAL  end1_cyc_dlyncs_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_gen_cntr_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_normal_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_reg_in_wire :	STD_LOGIC;
	 SIGNAL  end_add_cycle :	STD_LOGIC;
	 SIGNAL  end_add_cycle_mux_datab_wire :	STD_LOGIC;
	 SIGNAL  end_fast_read :	STD_LOGIC;
	 SIGNAL  end_one_cyc_pos :	STD_LOGIC;
	 SIGNAL  end_one_cycle :	STD_LOGIC;
	 SIGNAL  end_op_wire :	STD_LOGIC;
	 SIGNAL  end_operation :	STD_LOGIC;
	 SIGNAL  end_ophdly :	STD_LOGIC;
	 SIGNAL  end_pgwr_data :	STD_LOGIC;
	 SIGNAL  end_read :	STD_LOGIC;
	 SIGNAL  end_read_byte :	STD_LOGIC;
	 SIGNAL  end_wrstage :	STD_LOGIC;
	 SIGNAL  exb4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fast_read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fast_read_wire :	STD_LOGIC;
	 SIGNAL  freadwrv_sdoin :	STD_LOGIC;
	 SIGNAL  ill_erase_wire :	STD_LOGIC;
	 SIGNAL  ill_write_wire :	STD_LOGIC;
	 SIGNAL  illegal_erase_b4out_wire :	STD_LOGIC;
	 SIGNAL  illegal_write_b4out_wire :	STD_LOGIC;
	 SIGNAL  illegal_write_prot :	STD_LOGIC;
	 SIGNAL  in_operation :	STD_LOGIC;
	 SIGNAL  load_opcode :	STD_LOGIC;
	 SIGNAL  mask_prot :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mask_prot_add :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mask_prot_check :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mask_prot_comp_ntb :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mask_prot_comp_tb :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  memadd_sdoin :	STD_LOGIC;
	 SIGNAL  ncs_reg_ena_wire :	STD_LOGIC;
	 SIGNAL  not_busy :	STD_LOGIC;
	 SIGNAL  oe_wire :	STD_LOGIC;
	 SIGNAL  page_size_wire :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  pagewr_buf_not_empty :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  prot_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rden_wire :	STD_LOGIC;
	 SIGNAL  rdid_load :	STD_LOGIC;
	 SIGNAL  rdid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  reach_max_cnt :	STD_LOGIC;
	 SIGNAL  read_buf :	STD_LOGIC;
	 SIGNAL  read_bufdly :	STD_LOGIC;
	 SIGNAL  read_data_reg_in_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_rdid_wire :	STD_LOGIC;
	 SIGNAL  read_sid_wire :	STD_LOGIC;
	 SIGNAL  read_status_wire :	STD_LOGIC;
	 SIGNAL  read_wire :	STD_LOGIC;
	 SIGNAL  rflagstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rnvdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_sdoin :	STD_LOGIC;
	 SIGNAL  rstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  scein_wire :	STD_LOGIC;
	 SIGNAL  sdoin_wire :	STD_LOGIC;
	 SIGNAL  sec_erase_wire :	STD_LOGIC;
	 SIGNAL  sec_protect_wire :	STD_LOGIC;
	 SIGNAL  secprot_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  secprot_sdoin :	STD_LOGIC;
	 SIGNAL  serase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  shift_bytes_wire :	STD_LOGIC;
	 SIGNAL  shift_opcode :	STD_LOGIC;
	 SIGNAL  shift_opdata :	STD_LOGIC;
	 SIGNAL  shift_pgwr_data :	STD_LOGIC;
	 SIGNAL  st_busy_wire :	STD_LOGIC;
	 SIGNAL  stage2_wire :	STD_LOGIC;
	 SIGNAL  stage3_wire :	STD_LOGIC;
	 SIGNAL  stage4_wire :	STD_LOGIC;
	 SIGNAL  start_frpoll :	STD_LOGIC;
	 SIGNAL  start_poll :	STD_LOGIC;
	 SIGNAL  start_sppoll :	STD_LOGIC;
	 SIGNAL  start_wrpoll :	STD_LOGIC;
	 SIGNAL  to_sdoin_wire :	STD_LOGIC;
	 SIGNAL  wren_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wren_wire :	STD_LOGIC;
	 SIGNAL  write_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  write_prot_true :	STD_LOGIC;
	 SIGNAL  write_prot_true2 :	STD_LOGIC;
	 SIGNAL  write_sdoin :	STD_LOGIC;
	 SIGNAL  write_wire :	STD_LOGIC;
	 SIGNAL  wrvolatile_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_addr_range418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_range410w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range406w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range192w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range200w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_dataout_wire_range460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range205w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_exb4addr_opcode_range281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exb4addr_opcode_range187w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range245w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_range693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_add_range722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_check_range724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_ntb_range742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mask_prot_comp_tb_range744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_prot_wire_range679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range256w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range238w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range248w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range215w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range228w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range259w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range219w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range251w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range210w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range197w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range223w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range231w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 COMPONENT  a_graycounter
	 GENERIC 
	 (
		PVALUE	:	NATURAL := 0;
		WIDTH	:	NATURAL := 8;
		lpm_type	:	STRING := "a_graycounter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		q	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		qbin	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  scfifo
	 GENERIC 
	 (
		ADD_RAM_OUTPUT_REGISTER	:	STRING := "OFF";
		ALLOW_RWCYCLE_WHEN_FULL	:	STRING := "OFF";
		ALMOST_EMPTY_VALUE	:	NATURAL := 0;
		ALMOST_FULL_VALUE	:	NATURAL := 0;
		LPM_NUMWORDS	:	NATURAL;
		LPM_SHOWAHEAD	:	STRING := "OFF";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHU	:	NATURAL := 1;
		OVERFLOW_CHECKING	:	STRING := "ON";
		UNDERFLOW_CHECKING	:	STRING := "ON";
		USE_EAB	:	STRING := "ON";
		lpm_type	:	STRING := "scfifo"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		almost_empty	:	OUT STD_LOGIC;
		almost_full	:	OUT STD_LOGIC;
		clock	:	IN STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		empty	:	OUT STD_LOGIC;
		full	:	OUT STD_LOGIC;
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		rdreq	:	IN STD_LOGIC;
		sclr	:	IN STD_LOGIC := '0';
		usedw	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHU-1 DOWNTO 0);
		wrreq	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_w549w550w551w552w(0) <= wire_w_lg_w_lg_w549w550w551w(0) AND wire_w_lg_do_ex4baddr538w(0);
	wire_w_lg_w_lg_w549w550w551w(0) <= wire_w_lg_w549w550w(0) AND wire_w_lg_do_4baddr539w(0);
	wire_w_lg_w_lg_w799w800w801w(0) <= wire_w_lg_w799w800w(0) AND end_operation;
	wire_w_lg_w549w550w(0) <= wire_w549w(0) AND wire_w_lg_do_sec_prot540w(0);
	wire_w_lg_w799w800w(0) <= wire_w799w(0) AND wire_w_lg_do_ex4baddr538w(0);
	wire_w549w(0) <= wire_w_lg_w_lg_w_lg_w_lg_end_operation545w546w547w548w(0) AND wire_w_lg_do_bulk_erase541w(0);
	wire_w304w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode240w241w242w243w(0) AND wire_w_rdummyclk_opcode_range303w(0);
	loop0 : FOR i IN 0 TO 6 GENERATE 
		wire_w244w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode240w241w242w243w(0) AND wire_w_rdummyclk_opcode_range238w(i);
	END GENERATE loop0;
	wire_w302w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode233w234w235w236w(0) AND wire_w_wrvolatile_opcode_range301w(0);
	loop1 : FOR i IN 0 TO 6 GENERATE 
		wire_w237w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode233w234w235w236w(0) AND wire_w_wrvolatile_opcode_range231w(i);
	END GENERATE loop1;
	wire_w799w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write544w796w797w798w(0) AND wire_w_lg_do_4baddr539w(0);
	wire_w492w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read422w489w490w491w(0) AND end_read_byte;
	wire_w_lg_w_lg_w_lg_w_lg_end_operation545w546w547w548w(0) <= wire_w_lg_w_lg_w_lg_end_operation545w546w547w(0) AND wire_w_lg_do_die_erase542w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode201w202w203w288w(0) <= wire_w_lg_w_lg_w_lg_load_opcode201w202w203w(0) AND wire_w_berase_opcode_range287w(0);
	loop2 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode201w202w203w204w(i) <= wire_w_lg_w_lg_w_lg_load_opcode201w202w203w(0) AND wire_w_berase_opcode_range200w(i);
	END GENERATE loop2;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode206w207w208w290w(0) <= wire_w_lg_w_lg_w_lg_load_opcode206w207w208w(0) AND wire_w_derase_opcode_range289w(0);
	loop3 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode206w207w208w209w(i) <= wire_w_lg_w_lg_w_lg_load_opcode206w207w208w(0) AND wire_w_derase_opcode_range205w(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode240w241w242w243w(0) <= wire_w_lg_w_lg_w_lg_load_opcode240w241w242w(0) AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode211w212w213w292w(0) <= wire_w_lg_w_lg_w_lg_load_opcode211w212w213w(0) AND wire_w_serase_opcode_range291w(0);
	loop4 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode211w212w213w214w(i) <= wire_w_lg_w_lg_w_lg_load_opcode211w212w213w(0) AND wire_w_serase_opcode_range210w(i);
	END GENERATE loop4;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode252w253w254w310w(0) <= wire_w_lg_w_lg_w_lg_load_opcode252w253w254w(0) AND wire_w_secprot_opcode_range309w(0);
	loop5 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode252w253w254w255w(i) <= wire_w_lg_w_lg_w_lg_load_opcode252w253w254w(0) AND wire_w_secprot_opcode_range251w(i);
	END GENERATE loop5;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode233w234w235w236w(0) <= wire_w_lg_w_lg_w_lg_load_opcode233w234w235w(0) AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_read374w375w376w377w(0) <= wire_w_lg_w_lg_w_lg_do_read374w375w376w(0) AND end_one_cycle;
	wire_w_lg_w_lg_w_lg_w_lg_do_write544w796w797w798w(0) <= wire_w_lg_w_lg_w_lg_do_write544w796w797w(0) AND wire_w_lg_do_die_erase542w(0);
	wire_w_lg_w_lg_w_lg_w644w791w792w802w(0) <= wire_w_lg_w_lg_w644w791w792w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_w_lg_do_read422w489w490w491w(0) <= wire_w_lg_w_lg_w_lg_do_read422w489w490w(0) AND end_one_cyc_pos;
	wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase61w431w432w433w(0) <= wire_w_lg_w_lg_w_lg_do_sec_erase61w431w432w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_end_operation545w546w547w(0) <= wire_w_lg_w_lg_end_operation545w546w(0) AND wire_w_lg_do_sec_erase543w(0);
	wire_w_lg_w_lg_w_lg_load_opcode201w202w203w(0) <= wire_w_lg_w_lg_load_opcode201w202w(0) AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_w_lg_w_lg_load_opcode206w207w208w(0) <= wire_w_lg_w_lg_load_opcode206w207w(0) AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_w_lg_w_lg_load_opcode216w221w296w(0) <= wire_w_lg_w_lg_load_opcode216w221w(0) AND wire_w_rstat_opcode_range295w(0);
	loop6 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode216w221w222w(i) <= wire_w_lg_w_lg_load_opcode216w221w(0) AND wire_w_rstat_opcode_range219w(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_w_lg_load_opcode216w217w294w(0) <= wire_w_lg_w_lg_load_opcode216w217w(0) AND wire_w_rflagstat_opcode_range293w(0);
	loop7 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode216w217w218w(i) <= wire_w_lg_w_lg_load_opcode216w217w(0) AND wire_w_rflagstat_opcode_range215w(i);
	END GENERATE loop7;
	wire_w_lg_w_lg_w_lg_load_opcode240w241w242w(0) <= wire_w_lg_w_lg_load_opcode240w241w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_w_lg_load_opcode211w212w213w(0) <= wire_w_lg_w_lg_load_opcode211w212w(0) AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_w_lg_w_lg_load_opcode252w253w254w(0) <= wire_w_lg_w_lg_load_opcode252w253w(0) AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_w_lg_w_lg_load_opcode233w234w235w(0) <= wire_w_lg_w_lg_load_opcode233w234w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_w_lg_bp2_wire660w661w662w(0) <= wire_w_lg_w_lg_bp2_wire660w661w(0) AND wire_w_lg_bp0_wire658w(0);
	wire_w_lg_w_lg_w_lg_bp2_wire660w661w665w(0) <= wire_w_lg_w_lg_bp2_wire660w661w(0) AND bp0_wire;
	wire_w_lg_w_lg_w_lg_bp2_wire660w667w668w(0) <= wire_w_lg_w_lg_bp2_wire660w667w(0) AND wire_w_lg_bp0_wire658w(0);
	wire_w_lg_w_lg_w_lg_bp2_wire660w667w670w(0) <= wire_w_lg_w_lg_bp2_wire660w667w(0) AND bp0_wire;
	wire_w_lg_w_lg_w_lg_do_read374w375w376w(0) <= wire_w_lg_w_lg_do_read374w375w(0) AND wire_w_lg_w_lg_do_write70w372w(0);
	wire_w_lg_w_lg_w_lg_do_read374w375w434w(0) <= wire_w_lg_w_lg_do_read374w375w(0) AND clr_write_wire2;
	wire_w_lg_w_lg_w_lg_do_write544w796w797w(0) <= wire_w_lg_w_lg_do_write544w796w(0) AND wire_w_lg_do_bulk_erase541w(0);
	wire_w_lg_w_lg_w644w791w792w(0) <= wire_w_lg_w644w791w(0) AND wire_wrstage_cntr_w_lg_w_q_range636w637w(0);
	wire_w_lg_w_lg_w_lg_do_read422w489w490w(0) <= wire_w_lg_w_lg_do_read422w489w(0) AND wire_stage_cntr_w_lg_w_q_range108w113w(0);
	wire_w_lg_w_lg_w_lg_do_sec_erase61w431w432w(0) <= wire_w_lg_w_lg_do_sec_erase61w431w(0) AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_w_lg_bp2_wire672w673w(0) <= wire_w_lg_bp2_wire672w(0) AND wire_w_lg_bp0_wire658w(0);
	wire_w_lg_w_lg_bp2_wire672w675w(0) <= wire_w_lg_bp2_wire672w(0) AND bp0_wire;
	wire_w_lg_w_lg_bp2_wire677w678w(0) <= wire_w_lg_bp2_wire677w(0) AND wire_w_lg_bp0_wire658w(0);
	wire_w_lg_w_lg_bp2_wire677w680w(0) <= wire_w_lg_bp2_wire677w(0) AND bp0_wire;
	wire_w_lg_w_lg_do_4baddr193w194w(0) <= wire_w_lg_do_4baddr193w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_do_ex4baddr188w189w(0) <= wire_w_lg_do_ex4baddr188w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_do_polling558w559w(0) <= wire_w_lg_do_polling558w(0) AND stage3_dly_reg;
	wire_w_lg_w_lg_do_read_stat129w130w(0) <= wire_w_lg_do_read_stat129w(0) AND wire_w_lg_w_lg_w125w126w127w(0);
	wire_w_lg_w_lg_do_write224w225w(0) <= wire_w_lg_do_write224w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_do_write70w353w(0) <= wire_w_lg_do_write70w(0) AND end_pgwr_data;
	wire_w_lg_w_lg_end_operation545w546w(0) <= wire_w_lg_end_operation545w(0) AND wire_w_lg_do_write544w(0);
	wire_w_lg_w_lg_end_read_byte496w508w(0) <= wire_w_lg_end_read_byte496w(0) AND wire_w_lg_end_operation507w(0);
	wire_w_lg_w_lg_load_opcode195w284w(0) <= wire_w_lg_load_opcode195w(0) AND wire_w_b4addr_opcode_range283w(0);
	loop8 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode195w196w(i) <= wire_w_lg_load_opcode195w(0) AND wire_w_b4addr_opcode_range192w(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_load_opcode190w282w(0) <= wire_w_lg_load_opcode190w(0) AND wire_w_exb4addr_opcode_range281w(0);
	loop9 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode190w191w(i) <= wire_w_lg_load_opcode190w(0) AND wire_w_exb4addr_opcode_range187w(i);
	END GENERATE loop9;
	wire_w_lg_w_lg_load_opcode226w298w(0) <= wire_w_lg_load_opcode226w(0) AND wire_w_write_opcode_range297w(0);
	loop10 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode226w227w(i) <= wire_w_lg_load_opcode226w(0) AND wire_w_write_opcode_range223w(i);
	END GENERATE loop10;
	wire_w_lg_w_lg_load_opcode201w202w(0) <= wire_w_lg_load_opcode201w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_load_opcode206w207w(0) <= wire_w_lg_load_opcode206w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_load_opcode246w306w(0) <= wire_w_lg_load_opcode246w(0) AND wire_w_fast_read_opcode_range305w(0);
	loop11 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode246w247w(i) <= wire_w_lg_load_opcode246w(0) AND wire_w_fast_read_opcode_range245w(i);
	END GENERATE loop11;
	wire_w_lg_w_lg_load_opcode249w308w(0) <= wire_w_lg_load_opcode249w(0) AND wire_w_read_opcode_range307w(0);
	loop12 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode249w250w(i) <= wire_w_lg_load_opcode249w(0) AND wire_w_read_opcode_range248w(i);
	END GENERATE loop12;
	wire_w_lg_w_lg_load_opcode229w300w(0) <= wire_w_lg_load_opcode229w(0) AND wire_w_rnvdummyclk_opcode_range299w(0);
	loop13 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode229w230w(i) <= wire_w_lg_load_opcode229w(0) AND wire_w_rnvdummyclk_opcode_range228w(i);
	END GENERATE loop13;
	wire_w_lg_w_lg_load_opcode257w312w(0) <= wire_w_lg_load_opcode257w(0) AND wire_w_rdid_opcode_range311w(0);
	loop14 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode257w258w(i) <= wire_w_lg_load_opcode257w(0) AND wire_w_rdid_opcode_range256w(i);
	END GENERATE loop14;
	wire_w_lg_w_lg_load_opcode260w314w(0) <= wire_w_lg_load_opcode260w(0) AND wire_w_rsid_opcode_range313w(0);
	loop15 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode260w261w(i) <= wire_w_lg_load_opcode260w(0) AND wire_w_rsid_opcode_range259w(i);
	END GENERATE loop15;
	wire_w_lg_w_lg_load_opcode216w221w(0) <= wire_w_lg_load_opcode216w(0) AND wire_w_lg_do_polling220w(0);
	wire_w_lg_w_lg_load_opcode216w217w(0) <= wire_w_lg_load_opcode216w(0) AND do_polling;
	wire_w_lg_w_lg_load_opcode240w241w(0) <= wire_w_lg_load_opcode240w(0) AND wire_w_lg_do_write_volatile239w(0);
	wire_w_lg_w_lg_load_opcode211w212w(0) <= wire_w_lg_load_opcode211w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_load_opcode252w253w(0) <= wire_w_lg_load_opcode252w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_load_opcode198w286w(0) <= wire_w_lg_load_opcode198w(0) AND wire_w_wren_opcode_range285w(0);
	loop16 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode198w199w(i) <= wire_w_lg_load_opcode198w(0) AND wire_w_wren_opcode_range197w(i);
	END GENERATE loop16;
	wire_w_lg_w_lg_load_opcode233w234w(0) <= wire_w_lg_load_opcode233w(0) AND wire_w_lg_do_read_volatile232w(0);
	wire_w_lg_w_lg_reach_max_cnt626w627w(0) <= wire_w_lg_reach_max_cnt626w(0) AND wren_wire;
	wire_w_lg_w_lg_stage3_wire52w53w(0) <= wire_w_lg_stage3_wire52w(0) AND do_wait_dummyclk;
	wire_w_lg_w_lg_start_poll360w361w(0) <= wire_w_lg_start_poll360w(0) AND do_polling;
	wire_w_lg_w_lg_bp2_wire660w661w(0) <= wire_w_lg_bp2_wire660w(0) AND wire_w_lg_bp1_wire659w(0);
	wire_w_lg_w_lg_bp2_wire660w667w(0) <= wire_w_lg_bp2_wire660w(0) AND bp1_wire;
	wire_w_lg_w_lg_do_read374w375w(0) <= wire_w_lg_do_read374w(0) AND wire_w_lg_do_fast_read373w(0);
	wire_w_lg_w_lg_do_write544w796w(0) <= wire_w_lg_do_write544w(0) AND wire_w_lg_do_sec_erase543w(0);
	loop17 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_read_bufdly580w581w(i) <= wire_w_lg_read_bufdly580w(0) AND wire_pgwrbuf_dataout_w_q_range579w(i);
	END GENERATE loop17;
	wire_w_lg_w_lg_w631w632w633w(0) <= wire_w_lg_w631w632w(0) AND end_wrstage;
	wire_w_lg_w644w791w(0) <= wire_w644w(0) AND wire_wrstage_cntr_w_q_range638w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w630w(0) <= wire_w_lg_w_lg_w_lg_do_write79w122w123w(0) AND wire_w_lg_write_prot_true629w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w136w(0) <= wire_w_lg_w_lg_w_lg_do_write79w122w123w(0) AND write_prot_true;
	wire_w_lg_w_lg_w_lg_do_write79w80w423w(0) <= wire_w_lg_w_lg_do_write79w80w(0) AND do_memadd;
	wire_w_lg_w_lg_do_read422w489w(0) <= wire_w_lg_do_read422w(0) AND wire_stage_cntr_w_q_range109w(0);
	wire_w_lg_w_lg_do_read_rdid131w132w(0) <= wire_w_lg_do_read_rdid131w(0) AND end_op_wire;
	wire_w_lg_w_lg_do_sec_erase61w431w(0) <= wire_w_lg_do_sec_erase61w(0) AND wire_w_lg_do_wren60w(0);
	wire_w_lg_w_lg_end_operation560w561w(0) <= wire_w_lg_end_operation560w(0) AND do_read_stat;
	wire_w_lg_w_lg_rden_wire427w428w(0) <= wire_w_lg_rden_wire427w(0) AND not_busy;
	wire_w_lg_addr_overdie417w(0) <= addr_overdie AND wire_w_addr_reg_overdie_range416w(0);
	loop18 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_addr_overdie407w(i) <= addr_overdie AND wire_w_addr_reg_overdie_range406w(i);
	END GENERATE loop18;
	wire_w_lg_bp2_wire672w(0) <= bp2_wire AND wire_w_lg_bp1_wire659w(0);
	wire_w_lg_bp2_wire677w(0) <= bp2_wire AND bp1_wire;
	wire_w_lg_do_4baddr193w(0) <= do_4baddr AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_do_bulk_erase354w(0) <= do_bulk_erase AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_do_ex4baddr188w(0) <= do_ex4baddr AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_do_polling558w(0) <= do_polling AND end_one_cyc_pos;
	wire_w_lg_do_read_nonvolatile340w(0) <= do_read_nonvolatile AND wire_addbyte_cntr_w_q_range175w(0);
	wire_w_lg_do_read_stat129w(0) <= do_read_stat AND wire_w_lg_start_poll128w(0);
	wire_w_lg_do_write224w(0) <= do_write AND wire_w_lg_do_read_stat59w(0);
	wire_w_lg_do_write77w(0) <= do_write AND wire_w_lg_w_pagewr_buf_not_empty_range75w76w(0);
	wire_w_lg_do_write70w(0) <= do_write AND shift_pgwr_data;
	wire_w_lg_end_operation545w(0) <= end_operation AND do_read_stat;
	wire_w_lg_end_read_byte496w(0) <= end_read_byte AND end_one_cyc_pos;
	wire_w_lg_load_opcode195w(0) <= load_opcode AND wire_w_lg_w_lg_do_4baddr193w194w(0);
	wire_w_lg_load_opcode190w(0) <= load_opcode AND wire_w_lg_w_lg_do_ex4baddr188w189w(0);
	wire_w_lg_load_opcode226w(0) <= load_opcode AND wire_w_lg_w_lg_do_write224w225w(0);
	wire_w_lg_load_opcode201w(0) <= load_opcode AND do_bulk_erase;
	wire_w_lg_load_opcode206w(0) <= load_opcode AND do_die_erase;
	wire_w_lg_load_opcode246w(0) <= load_opcode AND do_fast_read;
	wire_w_lg_load_opcode249w(0) <= load_opcode AND do_read;
	wire_w_lg_load_opcode229w(0) <= load_opcode AND do_read_nonvolatile;
	wire_w_lg_load_opcode257w(0) <= load_opcode AND do_read_rdid;
	wire_w_lg_load_opcode260w(0) <= load_opcode AND do_read_sid;
	wire_w_lg_load_opcode216w(0) <= load_opcode AND do_read_stat;
	wire_w_lg_load_opcode240w(0) <= load_opcode AND do_read_volatile;
	wire_w_lg_load_opcode211w(0) <= load_opcode AND do_sec_erase;
	wire_w_lg_load_opcode252w(0) <= load_opcode AND do_sec_prot;
	wire_w_lg_load_opcode198w(0) <= load_opcode AND do_wren;
	wire_w_lg_load_opcode233w(0) <= load_opcode AND do_write_volatile;
	wire_w_lg_not_busy419w(0) <= not_busy AND wire_w_addr_range418w(0);
	loop19 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_not_busy411w(i) <= not_busy AND wire_w_addr_range410w(i);
	END GENERATE loop19;
	wire_w_lg_reach_max_cnt626w(0) <= reach_max_cnt AND shift_bytes_wire;
	wire_w_lg_read_bufdly588w(0) <= read_bufdly AND wire_scfifo3_w_q_range587w(0);
	loop20 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_read_bufdly583w(i) <= read_bufdly AND wire_scfifo3_w_q_range582w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_shift_opcode186w(i) <= shift_opcode AND wire_asmi_opcode_reg_w_q_range185w(i);
	END GENERATE loop21;
	wire_w_lg_stage3_wire425w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_w_lg_do_write79w80w423w424w(0);
	wire_w_lg_stage3_wire456w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_do_read_stat453w454w455w(0);
	wire_w_lg_stage3_wire62w(0) <= stage3_wire AND wire_w_lg_do_sec_erase61w(0);
	wire_w_lg_stage3_wire52w(0) <= stage3_wire AND do_fast_read;
	loop22 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_stage3_wire409w(i) <= stage3_wire AND wire_addr_reg_w_q_range408w(i);
	END GENERATE loop22;
	wire_w_lg_stage4_wire458w(0) <= stage4_wire AND wire_w_lg_w_lg_do_read422w457w(0);
	wire_w_lg_stage4_wire426w(0) <= stage4_wire AND addr_overdie;
	wire_w_lg_start_poll360w(0) <= start_poll AND do_read_stat;
	wire_w_lg_w_mask_prot_range682w695w(0) <= wire_w_mask_prot_range682w(0) AND wire_addr_reg_w_q_range694w(0);
	wire_w_lg_w_mask_prot_range685w702w(0) <= wire_w_mask_prot_range685w(0) AND wire_addr_reg_w_q_range701w(0);
	wire_w_lg_w_mask_prot_range687w707w(0) <= wire_w_mask_prot_range687w(0) AND wire_addr_reg_w_q_range706w(0);
	wire_w_lg_w_mask_prot_range689w712w(0) <= wire_w_mask_prot_range689w(0) AND wire_addr_reg_w_q_range711w(0);
	wire_w_lg_w_mask_prot_range691w717w(0) <= wire_w_mask_prot_range691w(0) AND wire_addr_reg_w_q_range716w(0);
	wire_w_lg_w_mask_prot_range693w721w(0) <= wire_w_mask_prot_range693w(0) AND wire_addr_reg_w_q_range439w(0);
	wire_w_lg_w_lg_do_write70w372w(0) <= NOT wire_w_lg_do_write70w(0);
	wire_w_lg_w_lg_w125w126w127w(0) <= NOT wire_w_lg_w125w126w(0);
	wire_w_lg_addr_overdie521w(0) <= NOT addr_overdie;
	wire_w_lg_bp0_wire658w(0) <= NOT bp0_wire;
	wire_w_lg_bp1_wire659w(0) <= NOT bp1_wire;
	wire_w_lg_bp2_wire660w(0) <= NOT bp2_wire;
	wire_w_lg_buf_empty765w(0) <= NOT buf_empty;
	wire_w_lg_busy_wire3w(0) <= NOT busy_wire;
	wire_w_lg_clkin_wire45w(0) <= NOT clkin_wire;
	wire_w_lg_do_4baddr539w(0) <= NOT do_4baddr;
	wire_w_lg_do_bulk_erase541w(0) <= NOT do_bulk_erase;
	wire_w_lg_do_die_erase542w(0) <= NOT do_die_erase;
	wire_w_lg_do_ex4baddr538w(0) <= NOT do_ex4baddr;
	wire_w_lg_do_fast_read373w(0) <= NOT do_fast_read;
	wire_w_lg_do_memadd440w(0) <= NOT do_memadd;
	wire_w_lg_do_polling220w(0) <= NOT do_polling;
	wire_w_lg_do_read374w(0) <= NOT do_read;
	wire_w_lg_do_read_rdid58w(0) <= NOT do_read_rdid;
	wire_w_lg_do_read_stat59w(0) <= NOT do_read_stat;
	wire_w_lg_do_read_volatile232w(0) <= NOT do_read_volatile;
	wire_w_lg_do_sec_erase543w(0) <= NOT do_sec_erase;
	wire_w_lg_do_sec_prot540w(0) <= NOT do_sec_prot;
	wire_w_lg_do_wren60w(0) <= NOT do_wren;
	wire_w_lg_do_write544w(0) <= NOT do_write;
	wire_w_lg_do_write_volatile239w(0) <= NOT do_write_volatile;
	wire_w_lg_end_add_cycle90w(0) <= NOT end_add_cycle;
	wire_w_lg_end_fast_read84w(0) <= NOT end_fast_read;
	wire_w_lg_end_operation507w(0) <= NOT end_operation;
	wire_w_lg_end_ophdly46w(0) <= NOT end_ophdly;
	wire_w_lg_end_pgwr_data69w(0) <= NOT end_pgwr_data;
	wire_w_lg_end_read87w(0) <= NOT end_read;
	wire_w_lg_rden_wire523w(0) <= NOT rden_wire;
	wire_w_lg_reach_max_cnt590w(0) <= NOT reach_max_cnt;
	wire_w_lg_read_bufdly580w(0) <= NOT read_bufdly;
	wire_w_lg_read_rdid_wire12w(0) <= NOT read_rdid_wire;
	wire_w_lg_read_sid_wire11w(0) <= NOT read_sid_wire;
	wire_w_lg_read_status_wire26w(0) <= NOT read_status_wire;
	wire_w_lg_sec_protect_wire10w(0) <= NOT sec_protect_wire;
	wire_w_lg_st_busy_wire133w(0) <= NOT st_busy_wire;
	wire_w_lg_start_poll128w(0) <= NOT start_poll;
	wire_w_lg_write_prot_true629w(0) <= NOT write_prot_true;
	wire_w_lg_write_wire20w(0) <= NOT write_wire;
	wire_w_lg_w_pagewr_buf_not_empty_range75w76w(0) <= NOT wire_w_pagewr_buf_not_empty_range75w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w644w791w792w802w803w(0) <= wire_w_lg_w_lg_w_lg_w644w791w792w802w(0) OR write_prot_true;
	wire_w_lg_w_lg_w_lg_load_opcode260w314w315w(0) <= wire_w_lg_w_lg_load_opcode260w314w(0) OR wire_w_lg_w_lg_load_opcode257w312w(0);
	loop23 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode260w261w262w(i) <= wire_w_lg_w_lg_load_opcode260w261w(i) OR wire_w_lg_w_lg_load_opcode257w258w(i);
	END GENERATE loop23;
	wire_w631w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w630w(0) OR do_4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_do_write79w80w423w424w(0) <= wire_w_lg_w_lg_w_lg_do_write79w80w423w(0) OR wire_w_lg_do_read422w(0);
	wire_w_lg_w_lg_w_lg_end_operation560w561w562w(0) <= wire_w_lg_w_lg_end_operation560w561w(0) OR clr_rstat_wire;
	wire_w_lg_w_lg_w_lg_rden_wire427w428w429w(0) <= wire_w_lg_w_lg_rden_wire427w428w(0) OR wire_w_lg_stage4_wire426w(0);
	wire_w_lg_w_lg_not_busy419w420w(0) <= wire_w_lg_not_busy419w(0) OR wire_w_lg_addr_overdie417w(0);
	loop24 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_not_busy411w412w(i) <= wire_w_lg_not_busy411w(i) OR wire_w_lg_stage3_wire409w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_read_bufdly583w584w(i) <= wire_w_lg_read_bufdly583w(i) OR wire_w_lg_w_lg_read_bufdly580w581w(i);
	END GENERATE loop25;
	wire_w_lg_w_lg_stage4_wire458w459w(0) <= wire_w_lg_stage4_wire458w(0) OR wire_w_lg_stage3_wire456w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode260w314w315w316w(0) <= wire_w_lg_w_lg_w_lg_load_opcode260w314w315w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode252w253w254w310w(0);
	loop26 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode260w261w262w263w(i) <= wire_w_lg_w_lg_w_lg_load_opcode260w261w262w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode252w253w254w255w(i);
	END GENERATE loop26;
	wire_w_lg_w631w632w(0) <= wire_w631w(0) OR do_ex4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_rden_wire427w428w429w430w(0) <= wire_w_lg_w_lg_w_lg_rden_wire427w428w429w(0) OR wire_w_lg_stage3_wire425w(0);
	loop27 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_w_lg_not_busy411w412w413w(i) <= wire_w_lg_w_lg_not_busy411w412w(i) OR wire_w_lg_addr_overdie407w(i);
	END GENERATE loop27;
	wire_w317w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode260w314w315w316w(0) OR wire_w_lg_w_lg_load_opcode249w308w(0);
	loop28 : FOR i IN 0 TO 6 GENERATE 
		wire_w264w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode260w261w262w263w(i) OR wire_w_lg_w_lg_load_opcode249w250w(i);
	END GENERATE loop28;
	wire_w_lg_w317w318w(0) <= wire_w317w(0) OR wire_w_lg_w_lg_load_opcode246w306w(0);
	loop29 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w264w265w(i) <= wire_w264w(i) OR wire_w_lg_w_lg_load_opcode246w247w(i);
	END GENERATE loop29;
	wire_w_lg_w_lg_w317w318w319w(0) <= wire_w_lg_w317w318w(0) OR wire_w304w(0);
	loop30 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w264w265w266w(i) <= wire_w_lg_w264w265w(i) OR wire_w244w(i);
	END GENERATE loop30;
	wire_w_lg_w_lg_w_lg_w317w318w319w320w(0) <= wire_w_lg_w_lg_w317w318w319w(0) OR wire_w302w(0);
	loop31 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w264w265w266w267w(i) <= wire_w_lg_w_lg_w264w265w266w(i) OR wire_w237w(i);
	END GENERATE loop31;
	wire_w_lg_w_lg_w_lg_w_lg_w317w318w319w320w321w(0) <= wire_w_lg_w_lg_w_lg_w317w318w319w320w(0) OR wire_w_lg_w_lg_load_opcode229w300w(0);
	loop32 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w264w265w266w267w268w(i) <= wire_w_lg_w_lg_w_lg_w264w265w266w267w(i) OR wire_w_lg_w_lg_load_opcode229w230w(i);
	END GENERATE loop32;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w317w318w319w320w321w322w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w317w318w319w320w321w(0) OR wire_w_lg_w_lg_load_opcode226w298w(0);
	loop33 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w264w265w266w267w268w269w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w264w265w266w267w268w(i) OR wire_w_lg_w_lg_load_opcode226w227w(i);
	END GENERATE loop33;
	wire_w323w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w317w318w319w320w321w322w(0) OR wire_w_lg_w_lg_w_lg_load_opcode216w221w296w(0);
	loop34 : FOR i IN 0 TO 6 GENERATE 
		wire_w270w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w264w265w266w267w268w269w(i) OR wire_w_lg_w_lg_w_lg_load_opcode216w221w222w(i);
	END GENERATE loop34;
	wire_w_lg_w323w324w(0) <= wire_w323w(0) OR wire_w_lg_w_lg_w_lg_load_opcode216w217w294w(0);
	loop35 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w270w271w(i) <= wire_w270w(i) OR wire_w_lg_w_lg_w_lg_load_opcode216w217w218w(i);
	END GENERATE loop35;
	wire_w_lg_w_lg_w323w324w325w(0) <= wire_w_lg_w323w324w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode211w212w213w292w(0);
	loop36 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w270w271w272w(i) <= wire_w_lg_w270w271w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode211w212w213w214w(i);
	END GENERATE loop36;
	wire_w_lg_w_lg_w_lg_w323w324w325w326w(0) <= wire_w_lg_w_lg_w323w324w325w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode206w207w208w290w(0);
	loop37 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w270w271w272w273w(i) <= wire_w_lg_w_lg_w270w271w272w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode206w207w208w209w(i);
	END GENERATE loop37;
	wire_w_lg_w_lg_w_lg_w_lg_w323w324w325w326w327w(0) <= wire_w_lg_w_lg_w_lg_w323w324w325w326w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode201w202w203w288w(0);
	loop38 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w270w271w272w273w274w(i) <= wire_w_lg_w_lg_w_lg_w270w271w272w273w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode201w202w203w204w(i);
	END GENERATE loop38;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w323w324w325w326w327w328w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w323w324w325w326w327w(0) OR wire_w_lg_w_lg_load_opcode198w286w(0);
	loop39 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w270w271w272w273w274w275w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w270w271w272w273w274w(i) OR wire_w_lg_w_lg_load_opcode198w199w(i);
	END GENERATE loop39;
	wire_w329w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w323w324w325w326w327w328w(0) OR wire_w_lg_w_lg_load_opcode195w284w(0);
	loop40 : FOR i IN 0 TO 6 GENERATE 
		wire_w276w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w270w271w272w273w274w275w(i) OR wire_w_lg_w_lg_load_opcode195w196w(i);
	END GENERATE loop40;
	wire_w_lg_w329w330w(0) <= wire_w329w(0) OR wire_w_lg_w_lg_load_opcode190w282w(0);
	loop41 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w276w277w(i) <= wire_w276w(i) OR wire_w_lg_w_lg_load_opcode190w191w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w276w277w278w(i) <= wire_w_lg_w276w277w(i) OR wire_w_lg_shift_opcode186w(i);
	END GENERATE loop42;
	wire_w_lg_w_lg_w168w169w170w(0) <= wire_w_lg_w168w169w(0) OR do_read_nonvolatile;
	wire_w_lg_w168w169w(0) <= wire_w168w(0) OR do_fast_read;
	wire_w_lg_w125w126w(0) <= wire_w125w(0) OR do_ex4baddr;
	wire_w168w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read_sid164w165w166w167w(0) OR do_read;
	wire_w644w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w643w(0) OR do_ex4baddr;
	wire_w125w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w124w(0) OR do_4baddr;
	wire_w_lg_w690w692w(0) <= wire_w690w(0) OR wire_w_prot_wire_range679w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_read422w443w444w445w(0) <= wire_w_lg_w_lg_w_lg_do_read422w443w444w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_w_lg_do_read_sid164w165w166w167w(0) <= wire_w_lg_w_lg_w_lg_do_read_sid164w165w166w(0) OR do_read_rdid;
	wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w643w(0) <= wire_w_lg_w_lg_w_lg_do_write79w122w123w(0) OR do_4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w124w(0) <= wire_w_lg_w_lg_w_lg_do_write79w122w123w(0) OR do_fread_epcq;
	wire_w690w(0) <= wire_w_lg_w_lg_w_lg_w_prot_wire_range666w684w686w688w(0) OR wire_w_prot_wire_range676w(0);
	wire_w_lg_w_lg_w_lg_bp3_wire653w654w655w(0) <= wire_w_lg_w_lg_bp3_wire653w654w(0) OR bp0_wire;
	wire_w_lg_w_lg_w_lg_do_read422w443w444w(0) <= wire_w_lg_w_lg_do_read422w443w(0) OR do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read_sid164w165w166w(0) <= wire_w_lg_w_lg_do_read_sid164w165w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_do_read_stat453w454w455w(0) <= wire_w_lg_w_lg_do_read_stat453w454w(0) OR do_read_nonvolatile;
	wire_w_lg_w_lg_w_lg_do_sec_erase646w647w648w(0) <= wire_w_lg_w_lg_do_sec_erase646w647w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_do_write79w122w123w(0) <= wire_w_lg_w_lg_do_write79w122w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_w_prot_wire_range666w684w686w688w(0) <= wire_w_lg_w_lg_w_prot_wire_range666w684w686w(0) OR wire_w_prot_wire_range674w(0);
	wire_w_lg_w_lg_bp3_wire653w654w(0) <= wire_w_lg_bp3_wire653w(0) OR bp1_wire;
	wire_w_lg_w_lg_do_read422w457w(0) <= wire_w_lg_do_read422w(0) OR do_read_sid;
	wire_w_lg_w_lg_do_read422w443w(0) <= wire_w_lg_do_read422w(0) OR do_write;
	wire_w_lg_w_lg_do_read_sid164w165w(0) <= wire_w_lg_do_read_sid164w(0) OR do_sec_erase;
	wire_w_lg_w_lg_do_read_stat453w454w(0) <= wire_w_lg_do_read_stat453w(0) OR do_read_volatile;
	wire_w_lg_w_lg_do_sec_erase646w647w(0) <= wire_w_lg_do_sec_erase646w(0) OR do_bulk_erase;
	wire_w_lg_w_lg_do_write79w122w(0) <= wire_w_lg_do_write79w(0) OR do_bulk_erase;
	wire_w_lg_w_lg_do_write79w80w(0) <= wire_w_lg_do_write79w(0) OR do_die_erase;
	wire_w_lg_w_lg_read_bufdly577w578w(0) <= wire_w_lg_read_bufdly577w(0) OR clr_write_wire;
	wire_w_lg_w_lg_w_prot_wire_range666w684w686w(0) <= wire_w_lg_w_prot_wire_range666w684w(0) OR wire_w_prot_wire_range671w(0);
	wire_w_lg_bp3_wire653w(0) <= bp3_wire OR bp2_wire;
	wire_w_lg_data0out_wire461w(0) <= data0out_wire OR wire_w_dataout_wire_range460w(0);
	wire_w_lg_do_4baddr356w(0) <= do_4baddr OR wire_w_lg_do_ex4baddr355w(0);
	wire_w_lg_do_ex4baddr355w(0) <= do_ex4baddr OR wire_w_lg_do_bulk_erase354w(0);
	wire_w_lg_do_read422w(0) <= do_read OR do_fast_read;
	wire_w_lg_do_read_rdid131w(0) <= do_read_rdid OR wire_w_lg_w_lg_do_read_stat129w130w(0);
	wire_w_lg_do_read_sid164w(0) <= do_read_sid OR do_write;
	wire_w_lg_do_read_stat453w(0) <= do_read_stat OR do_read_rdid;
	wire_w_lg_do_sec_erase61w(0) <= do_sec_erase OR do_die_erase;
	wire_w_lg_do_sec_erase646w(0) <= do_sec_erase OR do_write;
	wire_w_lg_do_wren357w(0) <= do_wren OR wire_w_lg_do_4baddr356w(0);
	wire_w_lg_do_write79w(0) <= do_write OR do_sec_erase;
	wire_w_lg_end_operation560w(0) <= end_operation OR wire_w_lg_w_lg_do_polling558w559w(0);
	wire_w_lg_load_opcode332w(0) <= load_opcode OR shift_opcode;
	wire_w_lg_rden_wire427w(0) <= rden_wire OR wren_wire;
	wire_w_lg_read_bufdly577w(0) <= read_bufdly OR shift_pgwr_data;
	wire_w_lg_w_mask_prot_add_range703w731w(0) <= wire_w_mask_prot_add_range703w(0) OR wire_w_mask_prot_comp_tb_range727w(0);
	wire_w_lg_w_mask_prot_add_range708w735w(0) <= wire_w_mask_prot_add_range708w(0) OR wire_w_mask_prot_comp_tb_range732w(0);
	wire_w_lg_w_mask_prot_add_range713w739w(0) <= wire_w_mask_prot_add_range713w(0) OR wire_w_mask_prot_comp_tb_range736w(0);
	wire_w_lg_w_mask_prot_add_range718w743w(0) <= wire_w_mask_prot_add_range718w(0) OR wire_w_mask_prot_comp_tb_range740w(0);
	wire_w_lg_w_mask_prot_add_range722w747w(0) <= wire_w_mask_prot_add_range722w(0) OR wire_w_mask_prot_comp_tb_range744w(0);
	wire_w_lg_w_mask_prot_check_range705w729w(0) <= wire_w_mask_prot_check_range705w(0) OR wire_w_mask_prot_comp_ntb_range725w(0);
	wire_w_lg_w_mask_prot_check_range710w733w(0) <= wire_w_mask_prot_check_range710w(0) OR wire_w_mask_prot_comp_ntb_range730w(0);
	wire_w_lg_w_mask_prot_check_range715w737w(0) <= wire_w_mask_prot_check_range715w(0) OR wire_w_mask_prot_comp_ntb_range734w(0);
	wire_w_lg_w_mask_prot_check_range720w741w(0) <= wire_w_mask_prot_check_range720w(0) OR wire_w_mask_prot_comp_ntb_range738w(0);
	wire_w_lg_w_mask_prot_check_range724w745w(0) <= wire_w_mask_prot_check_range724w(0) OR wire_w_mask_prot_comp_ntb_range742w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range595w598w(0) <= wire_w_pagewr_buf_not_empty_range595w(0) OR wire_pgwr_data_cntr_w_q_range597w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range599w601w(0) <= wire_w_pagewr_buf_not_empty_range599w(0) OR wire_pgwr_data_cntr_w_q_range600w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range602w604w(0) <= wire_w_pagewr_buf_not_empty_range602w(0) OR wire_pgwr_data_cntr_w_q_range603w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range605w607w(0) <= wire_w_pagewr_buf_not_empty_range605w(0) OR wire_pgwr_data_cntr_w_q_range606w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range608w610w(0) <= wire_w_pagewr_buf_not_empty_range608w(0) OR wire_pgwr_data_cntr_w_q_range609w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range611w613w(0) <= wire_w_pagewr_buf_not_empty_range611w(0) OR wire_pgwr_data_cntr_w_q_range612w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range614w616w(0) <= wire_w_pagewr_buf_not_empty_range614w(0) OR wire_pgwr_data_cntr_w_q_range615w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range617w619w(0) <= wire_w_pagewr_buf_not_empty_range617w(0) OR wire_pgwr_data_cntr_w_q_range618w(0);
	wire_w_lg_w_prot_wire_range666w684w(0) <= wire_w_prot_wire_range666w(0) OR wire_w_prot_wire_range669w(0);
	wire_w_lg_w_mask_prot_range682w698w(0) <= wire_w_mask_prot_range682w(0) XOR wire_w_mask_prot_add_range696w(0);
	wire_w_lg_w_mask_prot_range685w704w(0) <= wire_w_mask_prot_range685w(0) XOR wire_w_mask_prot_add_range703w(0);
	wire_w_lg_w_mask_prot_range687w709w(0) <= wire_w_mask_prot_range687w(0) XOR wire_w_mask_prot_add_range708w(0);
	wire_w_lg_w_mask_prot_range689w714w(0) <= wire_w_mask_prot_range689w(0) XOR wire_w_mask_prot_add_range713w(0);
	wire_w_lg_w_mask_prot_range691w719w(0) <= wire_w_mask_prot_range691w(0) XOR wire_w_mask_prot_add_range718w(0);
	wire_w_lg_w_mask_prot_range693w723w(0) <= wire_w_mask_prot_range693w(0) XOR wire_w_mask_prot_add_range722w(0);
	add_rollover <= add_rollover_reg;
	addr_overdie <= '0';
	addr_overdie_pos <= '0';
	addr_reg_overdie <= (OTHERS => '0');
	asmi_dataoe <= oe_wire;
	asmi_dclk <= clkin_wire;
	asmi_scein <= scein_wire;
	asmi_sdoin <= sdoin_wire;
	b4addr_opcode <= (OTHERS => '0');
	be_write_prot <= ((do_bulk_erase OR do_die_erase) AND wire_w_lg_w_lg_w_lg_bp3_wire653w654w655w(0));
	berase_opcode <= (OTHERS => '0');
	bp0_wire <= statreg_int(2);
	bp1_wire <= statreg_int(3);
	bp2_wire <= statreg_int(4);
	bp3_wire <= statreg_int(6);
	buf_empty <= buf_empty_reg;
	busy <= (busy_wire OR busy_delay_reg);
	busy_wire <= ((((((((((((((do_read_rdid OR do_read_sid) OR do_read) OR do_fast_read) OR do_write) OR do_sec_prot) OR do_read_stat) OR do_sec_erase) OR do_bulk_erase) OR do_die_erase) OR do_4baddr) OR do_read_volatile) OR do_fread_epcq) OR do_read_nonvolatile) OR do_ex4baddr);
	clkin_wire <= clkin;
	clr_addmsb_wire <= ((wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w114w435w436w(0) OR wire_w_lg_w_lg_w_lg_do_read374w375w434w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase61w431w432w433w(0));
	clr_endrbyte_wire <= ((((wire_w_lg_do_read422w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR clr_read_wire2);
	clr_rdid_wire <= clr_rdid_reg;
	clr_read_wire <= clr_read_reg;
	clr_read_wire2 <= clr_read_reg2;
	clr_rstat_wire <= clr_rstat_reg;
	clr_write_wire <= clr_write_reg;
	clr_write_wire2 <= clr_write_reg2;
	cnt_bfend_wire_in <= (wire_gen_cntr_w_lg_w_q_range119w120w(0) AND wire_gen_cntr_q(0));
	data0out_wire <= asmi_dataout;
	data_valid <= data_valid_wire;
	data_valid_wire <= dvalid_reg2;
	dataout <= ( read_data_reg(7 DOWNTO 0));
	dataout_wire <= ( "0000");
	derase_opcode <= (OTHERS => '0');
	do_4baddr <= '0';
	do_bulk_erase <= '0';
	do_die_erase <= '0';
	do_ex4baddr <= '0';
	do_fast_read <= (((wire_w_lg_read_rdid_wire12w(0) AND wire_w_lg_read_sid_wire11w(0)) AND wire_w_lg_sec_protect_wire10w(0)) AND fast_read_wire);
	do_fread_epcq <= '0';
	do_freadwrv_polling <= '0';
	do_memadd <= do_wrmemadd_reg;
	do_polling <= ((do_write_polling OR do_sprot_polling) OR do_freadwrv_polling);
	do_read <= '0';
	do_read_nonvolatile <= '0';
	do_read_rdid <= read_rdid_wire;
	do_read_sid <= '0';
	do_read_stat <= ((((((((wire_w_lg_read_rdid_wire12w(0) AND wire_w_lg_read_sid_wire11w(0)) AND wire_w_lg_sec_protect_wire10w(0)) AND (NOT (read_wire OR fast_read_wire))) AND wire_w_lg_write_wire20w(0)) AND read_status_wire) OR do_write_rstat) OR do_sprot_rstat) OR do_write_volatile_rstat);
	do_read_volatile <= '0';
	do_sec_erase <= ((((((wire_w_lg_read_rdid_wire12w(0) AND wire_w_lg_read_sid_wire11w(0)) AND wire_w_lg_sec_protect_wire10w(0)) AND (NOT (read_wire OR fast_read_wire))) AND wire_w_lg_write_wire20w(0)) AND wire_w_lg_read_status_wire26w(0)) AND sec_erase_wire);
	do_sec_prot <= '0';
	do_secprot_wren <= '0';
	do_sprot_polling <= '0';
	do_sprot_rstat <= '0';
	do_wait_dummyclk <= '0';
	do_wren <= ((do_write_wren OR do_secprot_wren) OR do_write_volatile_wren);
	do_write <= ((((wire_w_lg_read_rdid_wire12w(0) AND wire_w_lg_read_sid_wire11w(0)) AND wire_w_lg_sec_protect_wire10w(0)) AND (NOT (read_wire OR fast_read_wire))) AND write_wire);
	do_write_polling <= wire_w_lg_w_lg_w644w791w792w(0);
	do_write_rstat <= write_rstat_reg;
	do_write_volatile <= '0';
	do_write_volatile_rstat <= '0';
	do_write_volatile_wren <= '0';
	do_write_wren <= ((NOT wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0));
	dummy_read_buf <= maxcnt_shift_reg2;
	end1_cyc_dlyncs_in_wire <= (((((((((wire_stage_cntr_w_lg_w_lg_w_q_range108w113w139w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND (NOT wire_gen_cntr_q(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range108w113w139w140w141w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w136w(0)) OR wire_w_lg_do_write77w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire133w(0)));
	end1_cyc_gen_cntr_wire <= (wire_gen_cntr_w_lg_w_q_range119w120w(0) AND (NOT wire_gen_cntr_q(0)));
	end1_cyc_normal_in_wire <= ((((((((((wire_stage_cntr_w_lg_w_lg_w_q_range108w113w139w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range108w113w139w140w141w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w136w(0)) OR wire_w_lg_do_write77w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire133w(0))) OR wire_w_lg_w_lg_do_read_rdid131w132w(0));
	end1_cyc_reg_in_wire <= wire_mux211_dataout;
	end_add_cycle <= wire_mux212_dataout;
	end_add_cycle_mux_datab_wire <= (wire_addbyte_cntr_q(2) AND wire_addbyte_cntr_q(1));
	end_fast_read <= end_read_reg;
	end_one_cyc_pos <= end1_cyc_reg2;
	end_one_cycle <= end1_cyc_reg;
	end_op_wire <= (((((((((((wire_stage_cntr_w_lg_w_q_range109w114w(0) AND ((wire_w_lg_w_lg_w_lg_w_lg_do_read374w375w376w377w(0) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read))) OR (wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w112w369w370w(0) AND wire_w_lg_do_polling220w(0))) OR ((((((do_read_rdid AND end_one_cyc_pos) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) AND wire_addbyte_cntr_q(2)) AND wire_addbyte_cntr_q(1)) AND wire_addbyte_cntr_w_lg_w_q_range178w179w(0))) OR (wire_w_lg_w_lg_start_poll360w361w(0) AND wire_w_lg_st_busy_wire133w(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range109w110w111w358w359w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write79w122w123w136w(0)) OR wire_w_lg_w_lg_do_write70w353w(0)) OR wire_w_lg_do_write77w(0)) OR wire_stage_cntr_w352w(0)) OR wire_stage_cntr_w_lg_w347w348w(0)) OR (wire_stage_cntr_w_lg_w_lg_w_q_range109w112w342w(0) AND ((do_write_volatile OR do_read_volatile) OR wire_w_lg_do_read_nonvolatile340w(0))));
	end_operation <= end_op_reg;
	end_ophdly <= end_op_hdlyreg;
	end_pgwr_data <= end_pgwrop_reg;
	end_read <= end_read_reg;
	end_read_byte <= (end_rbyte_reg AND wire_w_lg_addr_overdie521w(0));
	end_wrstage <= end_operation;
	exb4addr_opcode <= (OTHERS => '0');
	fast_read_opcode <= "00001011";
	fast_read_wire <= fast_read_reg;
	freadwrv_sdoin <= '0';
	ill_erase_wire <= ill_erase_reg;
	ill_write_wire <= ill_write_reg;
	illegal_erase <= ill_erase_wire;
	illegal_erase_b4out_wire <= (((do_sec_erase OR do_bulk_erase) OR do_die_erase) AND write_prot_true);
	illegal_write <= ill_write_wire;
	illegal_write_b4out_wire <= (((do_write AND write_prot_true) OR (illegal_write_prot AND write_prot_true2)) OR wire_w_lg_do_write77w(0));
	illegal_write_prot <= illegal_write_prot_reg;
	in_operation <= busy_wire;
	load_opcode <= ((((wire_stage_cntr_w_lg_w_q_range109w110w(0) AND wire_stage_cntr_w_lg_w_q_range108w113w(0)) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_w_lg_w_q_range117w118w(0)) AND wire_gen_cntr_q(0));
	mask_prot <= ( wire_w_lg_w690w692w & wire_w690w & wire_w_lg_w_lg_w_lg_w_prot_wire_range666w684w686w688w & wire_w_lg_w_lg_w_prot_wire_range666w684w686w & wire_w_lg_w_prot_wire_range666w684w & prot_wire(1));
	mask_prot_add <= ( wire_w_lg_w_mask_prot_range693w721w & wire_w_lg_w_mask_prot_range691w717w & wire_w_lg_w_mask_prot_range689w712w & wire_w_lg_w_mask_prot_range687w707w & wire_w_lg_w_mask_prot_range685w702w & wire_w_lg_w_mask_prot_range682w695w);
	mask_prot_check <= ( wire_w_lg_w_mask_prot_range693w723w & wire_w_lg_w_mask_prot_range691w719w & wire_w_lg_w_mask_prot_range689w714w & wire_w_lg_w_mask_prot_range687w709w & wire_w_lg_w_mask_prot_range685w704w & wire_w_lg_w_mask_prot_range682w698w);
	mask_prot_comp_ntb <= ( wire_w_lg_w_mask_prot_check_range724w745w & wire_w_lg_w_mask_prot_check_range720w741w & wire_w_lg_w_mask_prot_check_range715w737w & wire_w_lg_w_mask_prot_check_range710w733w & wire_w_lg_w_mask_prot_check_range705w729w & mask_prot_check(0));
	mask_prot_comp_tb <= ( wire_w_lg_w_mask_prot_add_range722w747w & wire_w_lg_w_mask_prot_add_range718w743w & wire_w_lg_w_mask_prot_add_range713w739w & wire_w_lg_w_mask_prot_add_range708w735w & wire_w_lg_w_mask_prot_add_range703w731w & mask_prot_add(0));
	memadd_sdoin <= add_msb_reg;
	ncs_reg_ena_wire <= (((wire_stage_cntr_w_lg_w_lg_w_q_range109w110w111w(0) AND end_one_cyc_pos) OR addr_overdie_pos) OR end_operation);
	not_busy <= busy_det_reg;
	oe_wire <= '0';
	page_size_wire <= "100000000";
	pagewr_buf_not_empty <= ( wire_w_lg_w_pagewr_buf_not_empty_range617w619w & wire_w_lg_w_pagewr_buf_not_empty_range614w616w & wire_w_lg_w_pagewr_buf_not_empty_range611w613w & wire_w_lg_w_pagewr_buf_not_empty_range608w610w & wire_w_lg_w_pagewr_buf_not_empty_range605w607w & wire_w_lg_w_pagewr_buf_not_empty_range602w604w & wire_w_lg_w_pagewr_buf_not_empty_range599w601w & wire_w_lg_w_pagewr_buf_not_empty_range595w598w & wire_pgwr_data_cntr_q(0));
	prot_wire <= ( wire_w_lg_w_lg_bp2_wire677w680w & wire_w_lg_w_lg_bp2_wire677w678w & wire_w_lg_w_lg_bp2_wire672w675w & wire_w_lg_w_lg_bp2_wire672w673w & wire_w_lg_w_lg_w_lg_bp2_wire660w667w670w & wire_w_lg_w_lg_w_lg_bp2_wire660w667w668w & wire_w_lg_w_lg_w_lg_bp2_wire660w661w665w & wire_w_lg_w_lg_w_lg_bp2_wire660w661w662w);
	rden_wire <= rden;
	rdid_load <= (end_operation AND do_read_rdid);
	rdid_opcode <= "10011111";
	rdid_out <= ( rdid_out_reg(7 DOWNTO 0));
	rdummyclk_opcode <= (OTHERS => '0');
	reach_max_cnt <= max_cnt_reg;
	read_address <= ( read_add_reg(23 DOWNTO 0));
	read_buf <= (((((end_one_cycle AND do_write) AND wire_w_lg_do_read_stat59w(0)) AND wire_w_lg_do_wren60w(0)) AND (wire_stage_cntr_w_lg_w_q_range109w114w(0) OR wire_addbyte_cntr_w_lg_w_q_range175w180w(0))) AND wire_w_lg_buf_empty765w(0));
	read_bufdly <= read_bufdly_reg;
	read_data_reg_in_wire <= ( read_dout_reg(7 DOWNTO 0));
	read_opcode <= (OTHERS => '0');
	read_rdid_wire <= read_rdid_reg;
	read_sid_wire <= '0';
	read_status_wire <= read_status_reg;
	read_wire <= '0';
	rflagstat_opcode <= "00000101";
	rnvdummyclk_opcode <= (OTHERS => '0');
	rsid_opcode <= (OTHERS => '0');
	rsid_sdoin <= '0';
	rstat_opcode <= "00000101";
	scein_wire <= wire_ncs_reg_w_lg_q395w(0);
	sdoin_wire <= to_sdoin_wire;
	sec_erase_wire <= sec_erase_reg;
	sec_protect_wire <= '0';
	secprot_opcode <= (OTHERS => '0');
	secprot_sdoin <= '0';
	serase_opcode <= "11011000";
	shift_bytes_wire <= shift_bytes;
	shift_opcode <= shift_op_reg;
	shift_opdata <= stage2_wire;
	shift_pgwr_data <= shftpgwr_data_reg;
	st_busy_wire <= statreg_int(0);
	stage2_wire <= stage2_reg;
	stage3_wire <= stage3_reg;
	stage4_wire <= stage4_reg;
	start_frpoll <= '0';
	start_poll <= ((start_wrpoll OR start_sppoll) OR start_frpoll);
	start_sppoll <= '0';
	start_wrpoll <= start_wrpoll_reg2;
	status_out <= ( statreg_out(7 DOWNTO 0));
	to_sdoin_wire <= ((((((shift_opdata AND asmi_opcode_reg(7)) OR rsid_sdoin) OR memadd_sdoin) OR write_sdoin) OR secprot_sdoin) OR freadwrv_sdoin);
	wren_opcode <= "00000110";
	wren_wire <= '1';
	write_opcode <= "00000010";
	write_prot_true <= write_prot_reg;
	write_prot_true2 <= write_prot_reg2;
	write_sdoin <= ((((do_write AND stage4_wire) AND wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0)) AND pgwrbuf_dataout(7));
	write_wire <= write_reg;
	wrvolatile_opcode <= (OTHERS => '0');
	wire_w_addr_range418w(0) <= addr(0);
	wire_w_addr_range410w <= addr(23 DOWNTO 1);
	wire_w_addr_reg_overdie_range416w(0) <= addr_reg_overdie(0);
	wire_w_addr_reg_overdie_range406w <= addr_reg_overdie(23 DOWNTO 1);
	wire_w_b4addr_opcode_range283w(0) <= b4addr_opcode(0);
	wire_w_b4addr_opcode_range192w <= b4addr_opcode(7 DOWNTO 1);
	wire_w_berase_opcode_range287w(0) <= berase_opcode(0);
	wire_w_berase_opcode_range200w <= berase_opcode(7 DOWNTO 1);
	wire_w_dataout_wire_range460w(0) <= dataout_wire(1);
	wire_w_derase_opcode_range289w(0) <= derase_opcode(0);
	wire_w_derase_opcode_range205w <= derase_opcode(7 DOWNTO 1);
	wire_w_exb4addr_opcode_range281w(0) <= exb4addr_opcode(0);
	wire_w_exb4addr_opcode_range187w <= exb4addr_opcode(7 DOWNTO 1);
	wire_w_fast_read_opcode_range305w(0) <= fast_read_opcode(0);
	wire_w_fast_read_opcode_range245w <= fast_read_opcode(7 DOWNTO 1);
	wire_w_mask_prot_range682w(0) <= mask_prot(0);
	wire_w_mask_prot_range685w(0) <= mask_prot(1);
	wire_w_mask_prot_range687w(0) <= mask_prot(2);
	wire_w_mask_prot_range689w(0) <= mask_prot(3);
	wire_w_mask_prot_range691w(0) <= mask_prot(4);
	wire_w_mask_prot_range693w(0) <= mask_prot(5);
	wire_w_mask_prot_add_range696w(0) <= mask_prot_add(0);
	wire_w_mask_prot_add_range703w(0) <= mask_prot_add(1);
	wire_w_mask_prot_add_range708w(0) <= mask_prot_add(2);
	wire_w_mask_prot_add_range713w(0) <= mask_prot_add(3);
	wire_w_mask_prot_add_range718w(0) <= mask_prot_add(4);
	wire_w_mask_prot_add_range722w(0) <= mask_prot_add(5);
	wire_w_mask_prot_check_range705w(0) <= mask_prot_check(1);
	wire_w_mask_prot_check_range710w(0) <= mask_prot_check(2);
	wire_w_mask_prot_check_range715w(0) <= mask_prot_check(3);
	wire_w_mask_prot_check_range720w(0) <= mask_prot_check(4);
	wire_w_mask_prot_check_range724w(0) <= mask_prot_check(5);
	wire_w_mask_prot_comp_ntb_range725w(0) <= mask_prot_comp_ntb(0);
	wire_w_mask_prot_comp_ntb_range730w(0) <= mask_prot_comp_ntb(1);
	wire_w_mask_prot_comp_ntb_range734w(0) <= mask_prot_comp_ntb(2);
	wire_w_mask_prot_comp_ntb_range738w(0) <= mask_prot_comp_ntb(3);
	wire_w_mask_prot_comp_ntb_range742w(0) <= mask_prot_comp_ntb(4);
	wire_w_mask_prot_comp_tb_range727w(0) <= mask_prot_comp_tb(0);
	wire_w_mask_prot_comp_tb_range732w(0) <= mask_prot_comp_tb(1);
	wire_w_mask_prot_comp_tb_range736w(0) <= mask_prot_comp_tb(2);
	wire_w_mask_prot_comp_tb_range740w(0) <= mask_prot_comp_tb(3);
	wire_w_mask_prot_comp_tb_range744w(0) <= mask_prot_comp_tb(4);
	wire_w_pagewr_buf_not_empty_range595w(0) <= pagewr_buf_not_empty(0);
	wire_w_pagewr_buf_not_empty_range599w(0) <= pagewr_buf_not_empty(1);
	wire_w_pagewr_buf_not_empty_range602w(0) <= pagewr_buf_not_empty(2);
	wire_w_pagewr_buf_not_empty_range605w(0) <= pagewr_buf_not_empty(3);
	wire_w_pagewr_buf_not_empty_range608w(0) <= pagewr_buf_not_empty(4);
	wire_w_pagewr_buf_not_empty_range611w(0) <= pagewr_buf_not_empty(5);
	wire_w_pagewr_buf_not_empty_range614w(0) <= pagewr_buf_not_empty(6);
	wire_w_pagewr_buf_not_empty_range617w(0) <= pagewr_buf_not_empty(7);
	wire_w_pagewr_buf_not_empty_range75w(0) <= pagewr_buf_not_empty(8);
	wire_w_prot_wire_range666w(0) <= prot_wire(1);
	wire_w_prot_wire_range669w(0) <= prot_wire(2);
	wire_w_prot_wire_range671w(0) <= prot_wire(3);
	wire_w_prot_wire_range674w(0) <= prot_wire(4);
	wire_w_prot_wire_range676w(0) <= prot_wire(5);
	wire_w_prot_wire_range679w(0) <= prot_wire(6);
	wire_w_rdid_opcode_range311w(0) <= rdid_opcode(0);
	wire_w_rdid_opcode_range256w <= rdid_opcode(7 DOWNTO 1);
	wire_w_rdummyclk_opcode_range303w(0) <= rdummyclk_opcode(0);
	wire_w_rdummyclk_opcode_range238w <= rdummyclk_opcode(7 DOWNTO 1);
	wire_w_read_opcode_range307w(0) <= read_opcode(0);
	wire_w_read_opcode_range248w <= read_opcode(7 DOWNTO 1);
	wire_w_rflagstat_opcode_range293w(0) <= rflagstat_opcode(0);
	wire_w_rflagstat_opcode_range215w <= rflagstat_opcode(7 DOWNTO 1);
	wire_w_rnvdummyclk_opcode_range299w(0) <= rnvdummyclk_opcode(0);
	wire_w_rnvdummyclk_opcode_range228w <= rnvdummyclk_opcode(7 DOWNTO 1);
	wire_w_rsid_opcode_range313w(0) <= rsid_opcode(0);
	wire_w_rsid_opcode_range259w <= rsid_opcode(7 DOWNTO 1);
	wire_w_rstat_opcode_range295w(0) <= rstat_opcode(0);
	wire_w_rstat_opcode_range219w <= rstat_opcode(7 DOWNTO 1);
	wire_w_secprot_opcode_range309w(0) <= secprot_opcode(0);
	wire_w_secprot_opcode_range251w <= secprot_opcode(7 DOWNTO 1);
	wire_w_serase_opcode_range291w(0) <= serase_opcode(0);
	wire_w_serase_opcode_range210w <= serase_opcode(7 DOWNTO 1);
	wire_w_wren_opcode_range285w(0) <= wren_opcode(0);
	wire_w_wren_opcode_range197w <= wren_opcode(7 DOWNTO 1);
	wire_w_write_opcode_range297w(0) <= write_opcode(0);
	wire_w_write_opcode_range223w <= write_opcode(7 DOWNTO 1);
	wire_w_wrvolatile_opcode_range301w(0) <= wrvolatile_opcode(0);
	wire_w_wrvolatile_opcode_range231w <= wrvolatile_opcode(7 DOWNTO 1);
	wire_addbyte_cntr_w_lg_w_q_range175w180w(0) <= wire_addbyte_cntr_w_q_range175w(0) AND wire_addbyte_cntr_w_lg_w_q_range178w179w(0);
	wire_addbyte_cntr_w_lg_w_q_range178w179w(0) <= NOT wire_addbyte_cntr_w_q_range178w(0);
	wire_addbyte_cntr_clk_en <= wire_stage_cntr_w174w(0);
	wire_stage_cntr_w174w(0) <= ((wire_stage_cntr_w_lg_w_lg_w_q_range109w112w171w(0) AND wire_w_lg_w_lg_w168w169w170w(0)) OR addr_overdie) OR end_operation;
	wire_addbyte_cntr_clock <= wire_w_lg_clkin_wire45w(0);
	wire_addbyte_cntr_sclr <= wire_w_lg_end_operation107w(0);
	wire_w_lg_end_operation107w(0) <= end_operation OR addr_overdie;
	wire_addbyte_cntr_w_q_range178w(0) <= wire_addbyte_cntr_q(0);
	wire_addbyte_cntr_w_q_range175w(0) <= wire_addbyte_cntr_q(1);
	addbyte_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_addbyte_cntr_clk_en,
		clock => wire_addbyte_cntr_clock,
		q => wire_addbyte_cntr_q,
		sclr => wire_addbyte_cntr_sclr
	  );
	wire_gen_cntr_w_lg_w_q_range119w120w(0) <= wire_gen_cntr_w_q_range119w(0) AND wire_gen_cntr_w_lg_w_q_range117w118w(0);
	wire_gen_cntr_w_lg_w_q_range117w118w(0) <= NOT wire_gen_cntr_w_q_range117w(0);
	wire_gen_cntr_clk_en <= wire_w_lg_w_lg_w_lg_in_operation47w48w49w(0);
	wire_w_lg_w_lg_w_lg_in_operation47w48w49w(0) <= ((in_operation AND wire_w_lg_end_ophdly46w(0)) OR do_wait_dummyclk) OR addr_overdie;
	wire_gen_cntr_sclr <= wire_w_lg_w_lg_end1_cyc_reg_in_wire50w51w(0);
	wire_w_lg_w_lg_end1_cyc_reg_in_wire50w51w(0) <= (end1_cyc_reg_in_wire OR addr_overdie) OR do_wait_dummyclk;
	wire_gen_cntr_w_q_range117w(0) <= wire_gen_cntr_q(1);
	wire_gen_cntr_w_q_range119w(0) <= wire_gen_cntr_q(2);
	gen_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_gen_cntr_clk_en,
		clock => clkin_wire,
		q => wire_gen_cntr_q,
		sclr => wire_gen_cntr_sclr
	  );
	wire_stage_cntr_w_lg_w347w348w(0) <= wire_stage_cntr_w347w(0) AND end_one_cycle;
	wire_stage_cntr_w347w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range109w112w344w345w346w(0) AND end_add_cycle;
	wire_stage_cntr_w352w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range109w112w349w350w351w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range109w112w344w345w346w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w112w344w345w(0) AND wire_w_lg_do_read_stat59w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range109w112w349w350w351w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w112w349w350w(0) AND wire_w_lg_do_read_stat59w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range109w110w111w358w359w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w110w111w358w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w114w435w436w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range109w114w435w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w112w344w345w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range109w112w344w(0) AND wire_w_lg_do_wren60w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w112w369w370w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range109w112w369w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w112w349w350w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range109w112w349w(0) AND wire_w_lg_do_wren60w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range109w110w111w358w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range109w110w111w(0) AND wire_w_lg_do_wren357w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range109w114w435w(0) <= wire_stage_cntr_w_lg_w_q_range109w114w(0) AND end_add_cycle;
	wire_stage_cntr_w_lg_w_lg_w_q_range109w112w344w(0) <= wire_stage_cntr_w_lg_w_q_range109w112w(0) AND wire_w_lg_do_sec_erase61w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range109w112w369w(0) <= wire_stage_cntr_w_lg_w_q_range109w112w(0) AND do_read_stat;
	wire_stage_cntr_w_lg_w_lg_w_q_range109w112w349w(0) <= wire_stage_cntr_w_lg_w_q_range109w112w(0) AND do_sec_prot;
	wire_stage_cntr_w_lg_w_lg_w_q_range109w112w171w(0) <= wire_stage_cntr_w_lg_w_q_range109w112w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_q_range109w112w342w(0) <= wire_stage_cntr_w_lg_w_q_range109w112w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range108w113w139w140w141w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range108w113w139w140w(0) AND end1_cyc_gen_cntr_wire;
	wire_stage_cntr_w_lg_w_lg_w_q_range108w113w139w(0) <= wire_stage_cntr_w_lg_w_q_range108w113w(0) AND wire_stage_cntr_w_lg_w_q_range109w110w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range109w110w111w(0) <= wire_stage_cntr_w_lg_w_q_range109w110w(0) AND wire_stage_cntr_w_q_range108w(0);
	wire_stage_cntr_w_lg_w_q_range109w114w(0) <= wire_stage_cntr_w_q_range109w(0) AND wire_stage_cntr_w_lg_w_q_range108w113w(0);
	wire_stage_cntr_w_lg_w_q_range109w112w(0) <= wire_stage_cntr_w_q_range109w(0) AND wire_stage_cntr_w_q_range108w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range108w113w139w140w(0) <= NOT wire_stage_cntr_w_lg_w_lg_w_q_range108w113w139w(0);
	wire_stage_cntr_w_lg_w_q_range108w113w(0) <= NOT wire_stage_cntr_w_q_range108w(0);
	wire_stage_cntr_w_lg_w_q_range109w110w(0) <= NOT wire_stage_cntr_w_q_range109w(0);
	wire_stage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w103w104w105w106w(0);
	wire_w_lg_w_lg_w_lg_w103w104w105w106w(0) <= (((((((((((((in_operation AND end_one_cycle) AND (NOT (stage3_wire AND wire_w_lg_end_add_cycle90w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_read87w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_fast_read84w(0)))) AND (NOT ((wire_w_lg_w_lg_do_write79w80w(0) OR do_bulk_erase) AND write_prot_true))) AND (NOT wire_w_lg_do_write77w(0))) AND (NOT (stage3_wire AND st_busy_wire))) AND (NOT (wire_w_lg_do_write70w(0) AND wire_w_lg_end_pgwr_data69w(0)))) AND (NOT (stage2_wire AND do_wren))) AND (NOT (((wire_w_lg_stage3_wire62w(0) AND wire_w_lg_do_wren60w(0)) AND wire_w_lg_do_read_stat59w(0)) AND wire_w_lg_do_read_rdid58w(0)))) AND (NOT (stage3_wire AND ((do_write_volatile OR do_read_volatile) OR do_read_nonvolatile)))) OR wire_w_lg_w_lg_stage3_wire52w53w(0)) OR addr_overdie) OR end_ophdly;
	wire_stage_cntr_sclr <= wire_w_lg_end_operation107w(0);
	wire_stage_cntr_w_q_range108w(0) <= wire_stage_cntr_q(0);
	wire_stage_cntr_w_q_range109w(0) <= wire_stage_cntr_q(1);
	stage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_stage_cntr_clk_en,
		clock => clkin_wire,
		q => wire_stage_cntr_q,
		sclr => wire_stage_cntr_sclr
	  );
	wire_wrstage_cntr_w_lg_w_q_range638w639w(0) <= wire_wrstage_cntr_w_q_range638w(0) AND wire_wrstage_cntr_w_lg_w_q_range636w637w(0);
	wire_wrstage_cntr_w_lg_w_q_range636w637w(0) <= NOT wire_wrstage_cntr_w_q_range636w(0);
	wire_wrstage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w_lg_w631w632w633w634w635w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w631w632w633w634w635w(0) <= (wire_w_lg_w_lg_w631w632w633w(0) AND wire_w_lg_st_busy_wire133w(0)) OR clr_write_wire2;
	wire_wrstage_cntr_clock <= wire_w_lg_clkin_wire45w(0);
	wire_wrstage_cntr_w_q_range636w(0) <= wire_wrstage_cntr_q(0);
	wire_wrstage_cntr_w_q_range638w(0) <= wire_wrstage_cntr_q(1);
	wrstage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_wrstage_cntr_clk_en,
		clock => wire_wrstage_cntr_clock,
		q => wire_wrstage_cntr_q,
		sclr => clr_write_wire2
	  );
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN add_msb_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_add_msb_reg_ena = '1') THEN 
				IF (clr_addmsb_wire = '1') THEN add_msb_reg <= '0';
				ELSE add_msb_reg <= wire_addr_reg_w_q_range439w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_add_msb_reg_ena <= ((((wire_w_lg_w_lg_w_lg_w_lg_do_read422w443w444w445w(0) AND (NOT (wire_w_lg_w_lg_do_write79w80w(0) AND wire_w_lg_do_memadd440w(0)))) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) OR clr_addmsb_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN add_rollover_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN add_rollover_reg <= (wire_read_add_cntr_q(24) OR clr_read_wire2);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(0) = '1') THEN addr_reg(0) <= wire_addr_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(1) = '1') THEN addr_reg(1) <= wire_addr_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(2) = '1') THEN addr_reg(2) <= wire_addr_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(3) = '1') THEN addr_reg(3) <= wire_addr_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(4) = '1') THEN addr_reg(4) <= wire_addr_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(5) = '1') THEN addr_reg(5) <= wire_addr_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(6) = '1') THEN addr_reg(6) <= wire_addr_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(7) = '1') THEN addr_reg(7) <= wire_addr_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(8) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(8) = '1') THEN addr_reg(8) <= wire_addr_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(9) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(9) = '1') THEN addr_reg(9) <= wire_addr_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(10) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(10) = '1') THEN addr_reg(10) <= wire_addr_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(11) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(11) = '1') THEN addr_reg(11) <= wire_addr_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(12) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(12) = '1') THEN addr_reg(12) <= wire_addr_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(13) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(13) = '1') THEN addr_reg(13) <= wire_addr_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(14) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(14) = '1') THEN addr_reg(14) <= wire_addr_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(15) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(15) = '1') THEN addr_reg(15) <= wire_addr_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(16) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(16) = '1') THEN addr_reg(16) <= wire_addr_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(17) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(17) = '1') THEN addr_reg(17) <= wire_addr_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(18) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(18) = '1') THEN addr_reg(18) <= wire_addr_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(19) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(19) = '1') THEN addr_reg(19) <= wire_addr_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(20) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(20) = '1') THEN addr_reg(20) <= wire_addr_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(21) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(21) = '1') THEN addr_reg(21) <= wire_addr_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(22) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(22) = '1') THEN addr_reg(22) <= wire_addr_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(23) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(23) = '1') THEN addr_reg(23) <= wire_addr_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_addr_reg_d <= ( wire_w_lg_w_lg_w_lg_not_busy411w412w413w & wire_w_lg_w_lg_not_busy419w420w);
	loop43 : FOR i IN 0 TO 23 GENERATE
		wire_addr_reg_ena(i) <= wire_w_lg_w_lg_w_lg_w_lg_rden_wire427w428w429w430w(0);
	END GENERATE loop43;
	wire_addr_reg_w_q_range694w(0) <= addr_reg(18);
	wire_addr_reg_w_q_range701w(0) <= addr_reg(19);
	wire_addr_reg_w_q_range706w(0) <= addr_reg(20);
	wire_addr_reg_w_q_range711w(0) <= addr_reg(21);
	wire_addr_reg_w_q_range408w <= addr_reg(22 DOWNTO 0);
	wire_addr_reg_w_q_range716w(0) <= addr_reg(22);
	wire_addr_reg_w_q_range439w(0) <= addr_reg(23);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(0) = '1') THEN asmi_opcode_reg(0) <= wire_asmi_opcode_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(1) = '1') THEN asmi_opcode_reg(1) <= wire_asmi_opcode_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(2) = '1') THEN asmi_opcode_reg(2) <= wire_asmi_opcode_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(3) = '1') THEN asmi_opcode_reg(3) <= wire_asmi_opcode_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(4) = '1') THEN asmi_opcode_reg(4) <= wire_asmi_opcode_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(5) = '1') THEN asmi_opcode_reg(5) <= wire_asmi_opcode_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(6) = '1') THEN asmi_opcode_reg(6) <= wire_asmi_opcode_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(7) = '1') THEN asmi_opcode_reg(7) <= wire_asmi_opcode_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_asmi_opcode_reg_d <= ( wire_w_lg_w_lg_w276w277w278w & wire_w_lg_w329w330w);
	loop44 : FOR i IN 0 TO 7 GENERATE
		wire_asmi_opcode_reg_ena(i) <= wire_w_lg_load_opcode332w(0);
	END GENERATE loop44;
	wire_asmi_opcode_reg_w_q_range185w <= asmi_opcode_reg(6 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN buf_empty_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN buf_empty_reg <= wire_cmpr5_aeb;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN busy_delay_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (power_up_reg = '1') THEN busy_delay_reg <= busy_wire;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN busy_det_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN busy_det_reg <= wire_w_lg_busy_wire3w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_rdid_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rdid_reg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_read_reg <= ((do_read_sid OR do_sec_prot) OR end_operation);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN clr_read_reg2 <= clr_read_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_rstat_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN clr_rstat_reg <= ((end_operation OR do_read_sid) OR do_read);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_write_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_write_reg <= ((((((wire_w_lg_w_lg_w_lg_w_lg_w644w791w792w802w803w(0) OR wire_w_lg_do_write77w(0)) OR wire_w_lg_w_lg_w799w800w801w(0)) OR do_read_sid) OR do_sec_prot) OR do_read) OR do_fast_read);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_write_reg2 <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_write_reg2 <= clr_write_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN cnt_bfend_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN cnt_bfend_reg <= cnt_bfend_wire_in;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN do_wrmemadd_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN do_wrmemadd_reg <= (wire_wrstage_cntr_q(1) AND wire_wrstage_cntr_q(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_dvalid_reg_ena = '1') THEN 
				IF (wire_dvalid_reg_sclr = '1') THEN dvalid_reg <= '0';
				ELSE dvalid_reg <= wire_w_lg_end_read_byte496w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_dvalid_reg_ena <= wire_w_lg_do_read422w(0);
	wire_dvalid_reg_sclr <= (end_op_wire OR end_operation);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN dvalid_reg2 <= dvalid_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end1_cyc_reg <= end1_cyc_reg_in_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end1_cyc_reg2 <= end_one_cycle;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_hdlyreg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_op_hdlyreg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end_op_reg <= end_op_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_pgwrop_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_end_pgwrop_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN end_pgwrop_reg <= '0';
				ELSE end_pgwrop_reg <= buf_empty;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_end_pgwrop_reg_ena <= (((cnt_bfend_reg AND do_write) AND shift_pgwr_data) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_rbyte_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_end_rbyte_reg_ena = '1') THEN 
				IF (wire_end_rbyte_reg_sclr = '1') THEN end_rbyte_reg <= '0';
				ELSE end_rbyte_reg <= wire_w_lg_w_lg_w_lg_do_read422w489w490w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_end_rbyte_reg_ena <= ((wire_gen_cntr_w_lg_w_q_range119w120w(0) AND wire_gen_cntr_q(0)) OR clr_endrbyte_wire);
	wire_end_rbyte_reg_sclr <= (clr_endrbyte_wire OR addr_overdie);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_read_reg <= (((wire_w_lg_rden_wire523w(0) AND wire_w_lg_do_read422w(0)) AND data_valid_wire) AND end_read_byte);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN fast_read_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_fast_read_reg_ena = '1') THEN 
				IF (clr_read_wire = '1') THEN fast_read_reg <= '0';
				ELSE fast_read_reg <= fast_read;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_fast_read_reg_ena <= ((wire_w_lg_busy_wire3w(0) AND rden_wire) OR clr_read_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN ill_erase_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN ill_erase_reg <= (illegal_erase_dly_reg OR illegal_erase_b4out_wire);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN ill_write_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN ill_write_reg <= (illegal_write_dly_reg OR illegal_write_b4out_wire);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN illegal_erase_dly_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (power_up_reg = '1') THEN illegal_erase_dly_reg <= illegal_erase_b4out_wire;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN illegal_write_dly_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (power_up_reg = '1') THEN illegal_write_dly_reg <= illegal_write_b4out_wire;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN illegal_write_prot_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN illegal_write_prot_reg <= do_write;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN max_cnt_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN max_cnt_reg <= wire_cmpr4_aeb;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN maxcnt_shift_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN maxcnt_shift_reg <= (wire_w_lg_w_lg_reach_max_cnt626w627w(0) AND wire_w_lg_do_write544w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN maxcnt_shift_reg2 <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN maxcnt_shift_reg2 <= maxcnt_shift_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN ncs_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (ncs_reg_ena_wire = '1') THEN 
				IF (wire_ncs_reg_sclr = '1') THEN ncs_reg <= '0';
				ELSE ncs_reg <= '1';
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_ncs_reg_sclr <= (end_operation OR addr_overdie_pos);
	wire_ncs_reg_w_lg_q395w(0) <= NOT ncs_reg;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(0) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(0) <= '0';
				ELSE pgwrbuf_dataout(0) <= wire_pgwrbuf_dataout_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(1) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(1) <= '0';
				ELSE pgwrbuf_dataout(1) <= wire_pgwrbuf_dataout_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(2) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(2) <= '0';
				ELSE pgwrbuf_dataout(2) <= wire_pgwrbuf_dataout_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(3) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(3) <= '0';
				ELSE pgwrbuf_dataout(3) <= wire_pgwrbuf_dataout_d(3);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(4) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(4) <= '0';
				ELSE pgwrbuf_dataout(4) <= wire_pgwrbuf_dataout_d(4);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(5) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(5) <= '0';
				ELSE pgwrbuf_dataout(5) <= wire_pgwrbuf_dataout_d(5);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(6) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(6) <= '0';
				ELSE pgwrbuf_dataout(6) <= wire_pgwrbuf_dataout_d(6);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN pgwrbuf_dataout(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(7) = '1') THEN 
				IF (clr_write_wire = '1') THEN pgwrbuf_dataout(7) <= '0';
				ELSE pgwrbuf_dataout(7) <= wire_pgwrbuf_dataout_d(7);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_pgwrbuf_dataout_d <= ( wire_w_lg_w_lg_read_bufdly583w584w & wire_w_lg_read_bufdly588w);
	loop45 : FOR i IN 0 TO 7 GENERATE
		wire_pgwrbuf_dataout_ena(i) <= wire_w_lg_w_lg_read_bufdly577w578w(0);
	END GENERATE loop45;
	wire_pgwrbuf_dataout_w_q_range579w <= pgwrbuf_dataout(6 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN power_up_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN power_up_reg <= (busy_wire OR busy_delay_reg);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN rdid_out_reg <= (OTHERS => '0');
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (rdid_load = '1') THEN rdid_out_reg <= ( read_dout_reg(7 DOWNTO 0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(0) = '1') THEN read_add_reg(0) <= wire_read_add_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(1) = '1') THEN read_add_reg(1) <= wire_read_add_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(2) = '1') THEN read_add_reg(2) <= wire_read_add_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(3) = '1') THEN read_add_reg(3) <= wire_read_add_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(4) = '1') THEN read_add_reg(4) <= wire_read_add_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(5) = '1') THEN read_add_reg(5) <= wire_read_add_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(6) = '1') THEN read_add_reg(6) <= wire_read_add_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(7) = '1') THEN read_add_reg(7) <= wire_read_add_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(8) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(8) = '1') THEN read_add_reg(8) <= wire_read_add_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(9) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(9) = '1') THEN read_add_reg(9) <= wire_read_add_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(10) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(10) = '1') THEN read_add_reg(10) <= wire_read_add_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(11) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(11) = '1') THEN read_add_reg(11) <= wire_read_add_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(12) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(12) = '1') THEN read_add_reg(12) <= wire_read_add_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(13) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(13) = '1') THEN read_add_reg(13) <= wire_read_add_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(14) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(14) = '1') THEN read_add_reg(14) <= wire_read_add_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(15) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(15) = '1') THEN read_add_reg(15) <= wire_read_add_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(16) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(16) = '1') THEN read_add_reg(16) <= wire_read_add_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(17) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(17) = '1') THEN read_add_reg(17) <= wire_read_add_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(18) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(18) = '1') THEN read_add_reg(18) <= wire_read_add_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(19) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(19) = '1') THEN read_add_reg(19) <= wire_read_add_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(20) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(20) = '1') THEN read_add_reg(20) <= wire_read_add_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(21) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(21) = '1') THEN read_add_reg(21) <= wire_read_add_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(22) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(22) = '1') THEN read_add_reg(22) <= wire_read_add_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(23) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(23) = '1') THEN read_add_reg(23) <= wire_read_add_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_read_add_reg_d <= ( wire_read_add_cntr_q(23 DOWNTO 0));
	loop46 : FOR i IN 0 TO 23 GENERATE
		wire_read_add_reg_ena(i) <= wire_w_lg_w_lg_end_read_byte496w508w(0);
	END GENERATE loop46;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_bufdly_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN read_bufdly_reg <= read_buf;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(0) = '1') THEN read_data_reg(0) <= wire_read_data_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(1) = '1') THEN read_data_reg(1) <= wire_read_data_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(2) = '1') THEN read_data_reg(2) <= wire_read_data_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(3) = '1') THEN read_data_reg(3) <= wire_read_data_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(4) = '1') THEN read_data_reg(4) <= wire_read_data_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(5) = '1') THEN read_data_reg(5) <= wire_read_data_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(6) = '1') THEN read_data_reg(6) <= wire_read_data_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(7) = '1') THEN read_data_reg(7) <= wire_read_data_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_data_reg_d <= ( read_data_reg_in_wire(7 DOWNTO 0));
	loop47 : FOR i IN 0 TO 7 GENERATE
		wire_read_data_reg_ena(i) <= wire_w492w(0);
	END GENERATE loop47;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(0) = '1') THEN read_dout_reg(0) <= wire_read_dout_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(1) = '1') THEN read_dout_reg(1) <= wire_read_dout_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(2) = '1') THEN read_dout_reg(2) <= wire_read_dout_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(3) = '1') THEN read_dout_reg(3) <= wire_read_dout_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(4) = '1') THEN read_dout_reg(4) <= wire_read_dout_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(5) = '1') THEN read_dout_reg(5) <= wire_read_dout_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(6) = '1') THEN read_dout_reg(6) <= wire_read_dout_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(7) = '1') THEN read_dout_reg(7) <= wire_read_dout_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_dout_reg_d <= ( read_dout_reg(6 DOWNTO 0) & wire_w_lg_data0out_wire461w);
	loop48 : FOR i IN 0 TO 7 GENERATE
		wire_read_dout_reg_ena(i) <= wire_w_lg_w_lg_stage4_wire458w459w(0);
	END GENERATE loop48;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_rdid_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_rdid_reg_ena = '1') THEN 
				IF (clr_rdid_wire = '1') THEN read_rdid_reg <= '0';
				ELSE read_rdid_reg <= read_rdid;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_read_rdid_reg_ena <= (wire_w_lg_busy_wire3w(0) OR clr_rdid_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_status_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_status_reg_ena = '1') THEN 
				IF (clr_rstat_wire = '1') THEN read_status_reg <= '0';
				ELSE read_status_reg <= read_status;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_read_status_reg_ena <= (wire_w_lg_busy_wire3w(0) OR clr_rstat_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN sec_erase_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_sec_erase_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN sec_erase_reg <= '0';
				ELSE sec_erase_reg <= sector_erase;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_sec_erase_reg_ena <= ((wire_w_lg_busy_wire3w(0) AND wren_wire) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN shftpgwr_data_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
				IF (end_operation = '1') THEN shftpgwr_data_reg <= '0';
				ELSE shftpgwr_data_reg <= ((wire_stage_cntr_w_lg_w_q_range109w114w(0) AND wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0));
				END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN shift_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN shift_op_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range109w110w111w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage2_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage2_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range109w110w111w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage3_dly_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN stage3_dly_reg <= wire_stage_cntr_w_lg_w_q_range109w112w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage3_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage3_reg <= wire_stage_cntr_w_lg_w_q_range109w112w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage4_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage4_reg <= wire_stage_cntr_w_lg_w_q_range109w114w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN start_wrpoll_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_start_wrpoll_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN start_wrpoll_reg <= '0';
				ELSE start_wrpoll_reg <= wire_stage_cntr_w_lg_w_q_range109w112w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_start_wrpoll_reg_ena <= (((do_write_rstat AND do_polling) AND end_one_cycle) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN start_wrpoll_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
				IF (clr_write_wire = '1') THEN start_wrpoll_reg2 <= '0';
				ELSE start_wrpoll_reg2 <= start_wrpoll_reg;
				END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(0) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(0) <= '0';
				ELSE statreg_int(0) <= wire_statreg_int_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(1) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(1) <= '0';
				ELSE statreg_int(1) <= wire_statreg_int_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(2) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(2) <= '0';
				ELSE statreg_int(2) <= wire_statreg_int_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(3) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(3) <= '0';
				ELSE statreg_int(3) <= wire_statreg_int_d(3);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(4) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(4) <= '0';
				ELSE statreg_int(4) <= wire_statreg_int_d(4);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(5) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(5) <= '0';
				ELSE statreg_int(5) <= wire_statreg_int_d(5);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(6) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(6) <= '0';
				ELSE statreg_int(6) <= wire_statreg_int_d(6);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_int(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(7) = '1') THEN 
				IF (clr_rstat_wire = '1') THEN statreg_int(7) <= '0';
				ELSE statreg_int(7) <= wire_statreg_int_d(7);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_statreg_int_d <= ( read_dout_reg(7 DOWNTO 0));
	loop49 : FOR i IN 0 TO 7 GENERATE
		wire_statreg_int_ena(i) <= wire_w_lg_w_lg_w_lg_end_operation560w561w562w(0);
	END GENERATE loop49;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(0) = '1') THEN statreg_out(0) <= wire_statreg_out_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(1) = '1') THEN statreg_out(1) <= wire_statreg_out_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(2) = '1') THEN statreg_out(2) <= wire_statreg_out_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(3) = '1') THEN statreg_out(3) <= wire_statreg_out_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(4) = '1') THEN statreg_out(4) <= wire_statreg_out_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(5) = '1') THEN statreg_out(5) <= wire_statreg_out_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(6) = '1') THEN statreg_out(6) <= wire_statreg_out_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN statreg_out(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(7) = '1') THEN statreg_out(7) <= wire_statreg_out_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_statreg_out_d <= ( read_dout_reg(7 DOWNTO 0));
	loop50 : FOR i IN 0 TO 7 GENERATE
		wire_statreg_out_ena(i) <= wire_w_lg_w_lg_w_lg_w549w550w551w552w(0);
	END GENERATE loop50;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN write_prot_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_write_prot_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN write_prot_reg <= '0';
				ELSE write_prot_reg <= (((wire_w_lg_do_write79w(0) AND (NOT mask_prot_comp_ntb(5))) AND (NOT prot_wire(0))) OR be_write_prot);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_write_prot_reg_ena <= ((((wire_w_lg_w_lg_w_lg_do_sec_erase646w647w648w(0) AND (NOT wire_wrstage_cntr_q(1))) AND wire_wrstage_cntr_q(0)) AND end_ophdly) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN write_prot_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN write_prot_reg2 <= write_prot_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN write_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_write_reg_ena = '1') THEN 
				IF (clr_write_wire = '1') THEN write_reg <= '0';
				ELSE write_reg <= write;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_write_reg_ena <= ((wire_w_lg_busy_wire3w(0) AND wren_wire) OR clr_write_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN write_rstat_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
				IF (clr_write_wire = '1') THEN write_rstat_reg <= '0';
				ELSE write_rstat_reg <= (wire_w644w(0) AND (((NOT wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_w_lg_w_q_range636w637w(0)) OR wire_wrstage_cntr_w_lg_w_q_range638w639w(0)));
				END IF;
		END IF;
	END PROCESS;
	wire_cmpr4_dataa <= ( page_size_wire(8 DOWNTO 0));
	wire_cmpr4_datab <= ( wire_pgwr_data_cntr_q(8 DOWNTO 0));
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aeb => wire_cmpr4_aeb,
		dataa => wire_cmpr4_dataa,
		datab => wire_cmpr4_datab
	  );
	wire_cmpr5_dataa <= ( wire_pgwr_data_cntr_q(8 DOWNTO 0));
	wire_cmpr5_datab <= ( wire_pgwr_read_cntr_q(8 DOWNTO 0));
	cmpr5 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aeb => wire_cmpr5_aeb,
		dataa => wire_cmpr5_dataa,
		datab => wire_cmpr5_datab
	  );
	wire_pgwr_data_cntr_clk_en <= wire_w593w(0);
	wire_w593w(0) <= (((shift_bytes_wire AND wren_wire) AND wire_w_lg_reach_max_cnt590w(0)) AND wire_w_lg_do_write544w(0)) OR clr_write_wire2;
	wire_pgwr_data_cntr_w_q_range597w(0) <= wire_pgwr_data_cntr_q(1);
	wire_pgwr_data_cntr_w_q_range600w(0) <= wire_pgwr_data_cntr_q(2);
	wire_pgwr_data_cntr_w_q_range603w(0) <= wire_pgwr_data_cntr_q(3);
	wire_pgwr_data_cntr_w_q_range606w(0) <= wire_pgwr_data_cntr_q(4);
	wire_pgwr_data_cntr_w_q_range609w(0) <= wire_pgwr_data_cntr_q(5);
	wire_pgwr_data_cntr_w_q_range612w(0) <= wire_pgwr_data_cntr_q(6);
	wire_pgwr_data_cntr_w_q_range615w(0) <= wire_pgwr_data_cntr_q(7);
	wire_pgwr_data_cntr_w_q_range618w(0) <= wire_pgwr_data_cntr_q(8);
	pgwr_data_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 9
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_pgwr_data_cntr_clk_en,
		clock => clkin_wire,
		q => wire_pgwr_data_cntr_q,
		sclr => clr_write_wire2
	  );
	wire_pgwr_read_cntr_clk_en <= wire_w_lg_read_buf774w(0);
	wire_w_lg_read_buf774w(0) <= read_buf OR clr_write_wire2;
	pgwr_read_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 9
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_pgwr_read_cntr_clk_en,
		clock => clkin_wire,
		q => wire_pgwr_read_cntr_q,
		sclr => clr_write_wire2
	  );
	wire_read_add_cntr_clk_en <= wire_w_lg_w_lg_w_lg_rden_wire498w499w500w(0);
	wire_w_lg_w_lg_w_lg_rden_wire498w499w500w(0) <= ((rden_wire AND not_busy) OR data_valid_wire) OR add_rollover;
	wire_read_add_cntr_data <= ( "0" & addr(23 DOWNTO 0));
	wire_read_add_cntr_sload <= wire_w_lg_rden_wire498w(0);
	wire_w_lg_rden_wire498w(0) <= rden_wire AND not_busy;
	read_add_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 25
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_read_add_cntr_clk_en,
		clock => clkin_wire,
		data => wire_read_add_cntr_data,
		q => wire_read_add_cntr_q,
		sclr => add_rollover,
		sload => wire_read_add_cntr_sload
	  );
	wire_mux211_dataout <= end1_cyc_dlyncs_in_wire WHEN ((((do_write OR do_sec_prot) OR do_sec_erase) OR do_bulk_erase) OR do_die_erase) = '1'  ELSE end1_cyc_normal_in_wire;
	wire_mux212_dataout <= end_add_cycle_mux_datab_wire WHEN do_fast_read = '1'  ELSE wire_addbyte_cntr_w_lg_w_q_range175w180w(0);
	wire_scfifo3_data <= ( datain(7 DOWNTO 0));
	wire_scfifo3_rdreq <= wire_w_lg_read_buf576w(0);
	wire_w_lg_read_buf576w(0) <= read_buf OR dummy_read_buf;
	wire_scfifo3_wrreq <= wire_w_lg_w_lg_shift_bytes_wire574w575w(0);
	wire_w_lg_w_lg_shift_bytes_wire574w575w(0) <= (shift_bytes_wire AND wren_wire) AND wire_w_lg_do_write544w(0);
	wire_scfifo3_w_q_range582w <= wire_scfifo3_q(7 DOWNTO 1);
	wire_scfifo3_w_q_range587w(0) <= wire_scfifo3_q(0);
	scfifo3 :  scfifo
	  GENERIC MAP (
		LPM_NUMWORDS => 258,
		LPM_WIDTH => 8,
		LPM_WIDTHU => 9,
		USE_EAB => "ON"
	  )
	  PORT MAP ( 
		aclr => reset,
		clock => clkin_wire,
		data => wire_scfifo3_data,
		q => wire_scfifo3_q,
		rdreq => wire_scfifo3_rdreq,
		sclr => clr_write_wire2,
		wrreq => wire_scfifo3_wrreq
	  );

 END RTL; --altasmi_altasmi_parallel_pu03
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altasmi IS
	PORT
	(
		addr		: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		asmi_dataout		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		clkin		: IN STD_LOGIC ;
		datain		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		fast_read		: IN STD_LOGIC ;
		rden		: IN STD_LOGIC ;
		read_rdid		: IN STD_LOGIC ;
		read_status		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		sector_erase		: IN STD_LOGIC ;
		shift_bytes		: IN STD_LOGIC ;
		write		: IN STD_LOGIC ;
		asmi_dataoe		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		asmi_dclk		: OUT STD_LOGIC ;
		asmi_scein		: OUT STD_LOGIC ;
		asmi_sdoin		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		busy		: OUT STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		illegal_erase		: OUT STD_LOGIC ;
		illegal_write		: OUT STD_LOGIC ;
		rdid_out		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		read_address		: OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
		status_out		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END altasmi;


ARCHITECTURE RTL OF altasmi IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "ALTASMI_PARALLEL";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "data_width=STANDARD;epcs_type=EPCS128;intended_device_family=Arria II GX;lpm_hint=UNUSED;lpm_type=altasmi_parallel;page_size=256;port_bulk_erase=PORT_UNUSED;port_die_erase=PORT_UNUSED;port_en4b_addr=PORT_UNUSED;port_ex4b_addr=PORT_UNUSED;port_fast_read=PORT_USED;port_illegal_erase=PORT_USED;port_illegal_write=PORT_USED;port_rdid_out=PORT_USED;port_read_address=PORT_USED;port_read_dummyclk=PORT_UNUSED;port_read_rdid=PORT_USED;port_read_sid=PORT_UNUSED;port_read_status=PORT_USED;port_sector_erase=PORT_USED;port_sector_protect=PORT_UNUSED;port_shift_bytes=PORT_USED;port_wren=PORT_UNUSED;port_write=PORT_USED;use_asmiblock=OFF;use_eab=ON;write_dummy_clk=0;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (23 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC ;
	SIGNAL sub_wire8	: STD_LOGIC ;
	SIGNAL sub_wire9	: STD_LOGIC ;
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC ;



	COMPONENT altasmi_altasmi_parallel_pu03
	PORT (
			clkin	: IN STD_LOGIC ;
			data_valid	: OUT STD_LOGIC ;
			datain	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			fast_read	: IN STD_LOGIC ;
			illegal_erase	: OUT STD_LOGIC ;
			rden	: IN STD_LOGIC ;
			read_address	: OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
			asmi_sdoin	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			rdid_out	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			read_rdid	: IN STD_LOGIC ;
			addr	: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
			asmi_dataoe	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			asmi_dataout	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			asmi_dclk	: OUT STD_LOGIC ;
			asmi_scein	: OUT STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			read_status	: IN STD_LOGIC ;
			reset	: IN STD_LOGIC ;
			sector_erase	: IN STD_LOGIC ;
			status_out	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			write	: IN STD_LOGIC ;
			illegal_write	: OUT STD_LOGIC ;
			shift_bytes	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	data_valid    <= sub_wire0;
	illegal_erase    <= sub_wire1;
	read_address    <= sub_wire2(23 DOWNTO 0);
	asmi_sdoin    <= sub_wire3(0 DOWNTO 0);
	dataout    <= sub_wire4(7 DOWNTO 0);
	rdid_out    <= sub_wire5(7 DOWNTO 0);
	asmi_dataoe    <= sub_wire6(0 DOWNTO 0);
	asmi_dclk    <= sub_wire7;
	asmi_scein    <= sub_wire8;
	busy    <= sub_wire9;
	status_out    <= sub_wire10(7 DOWNTO 0);
	illegal_write    <= sub_wire11;

	altasmi_altasmi_parallel_pu03_component : altasmi_altasmi_parallel_pu03
	PORT MAP (
		clkin => clkin,
		datain => datain,
		fast_read => fast_read,
		rden => rden,
		read_rdid => read_rdid,
		addr => addr,
		asmi_dataout => asmi_dataout,
		read_status => read_status,
		reset => reset,
		sector_erase => sector_erase,
		write => write,
		shift_bytes => shift_bytes,
		data_valid => sub_wire0,
		illegal_erase => sub_wire1,
		read_address => sub_wire2,
		asmi_sdoin => sub_wire3,
		dataout => sub_wire4,
		rdid_out => sub_wire5,
		asmi_dataoe => sub_wire6,
		asmi_dclk => sub_wire7,
		asmi_scein => sub_wire8,
		busy => sub_wire9,
		status_out => sub_wire10,
		illegal_write => sub_wire11
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: CONSTANT: DATA_WIDTH STRING "STANDARD"
-- Retrieval info: CONSTANT: EPCS_TYPE STRING "EPCS128"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altasmi_parallel"
-- Retrieval info: CONSTANT: PAGE_SIZE NUMERIC "256"
-- Retrieval info: CONSTANT: PORT_BULK_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_DIE_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_EN4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_EX4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_FAST_READ STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_ERASE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_WRITE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_RDID_OUT STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_ADDRESS STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_DUMMYCLK STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_RDID STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_SID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_STATUS STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_SECTOR_ERASE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_SECTOR_PROTECT STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SHIFT_BYTES STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_WREN STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_WRITE STRING "PORT_USED"
-- Retrieval info: CONSTANT: USE_ASMIBLOCK STRING "OFF"
-- Retrieval info: CONSTANT: USE_EAB STRING "ON"
-- Retrieval info: CONSTANT: WRITE_DUMMY_CLK NUMERIC "0"
-- Retrieval info: USED_PORT: addr 0 0 24 0 INPUT NODEFVAL "addr[23..0]"
-- Retrieval info: CONNECT: @addr 0 0 24 0 addr 0 0 24 0
-- Retrieval info: USED_PORT: asmi_dataoe 0 0 1 0 OUTPUT NODEFVAL "asmi_dataoe[0..0]"
-- Retrieval info: CONNECT: asmi_dataoe 0 0 1 0 @asmi_dataoe 0 0 1 0
-- Retrieval info: USED_PORT: asmi_dataout 0 0 1 0 INPUT NODEFVAL "asmi_dataout[0..0]"
-- Retrieval info: CONNECT: @asmi_dataout 0 0 1 0 asmi_dataout 0 0 1 0
-- Retrieval info: USED_PORT: asmi_dclk 0 0 0 0 OUTPUT NODEFVAL "asmi_dclk"
-- Retrieval info: CONNECT: asmi_dclk 0 0 0 0 @asmi_dclk 0 0 0 0
-- Retrieval info: USED_PORT: asmi_scein 0 0 0 0 OUTPUT NODEFVAL "asmi_scein"
-- Retrieval info: CONNECT: asmi_scein 0 0 0 0 @asmi_scein 0 0 0 0
-- Retrieval info: USED_PORT: asmi_sdoin 0 0 1 0 OUTPUT NODEFVAL "asmi_sdoin[0..0]"
-- Retrieval info: CONNECT: asmi_sdoin 0 0 1 0 @asmi_sdoin 0 0 1 0
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: USED_PORT: clkin 0 0 0 0 INPUT NODEFVAL "clkin"
-- Retrieval info: CONNECT: @clkin 0 0 0 0 clkin 0 0 0 0
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: USED_PORT: datain 0 0 8 0 INPUT NODEFVAL "datain[7..0]"
-- Retrieval info: CONNECT: @datain 0 0 8 0 datain 0 0 8 0
-- Retrieval info: USED_PORT: dataout 0 0 8 0 OUTPUT NODEFVAL "dataout[7..0]"
-- Retrieval info: CONNECT: dataout 0 0 8 0 @dataout 0 0 8 0
-- Retrieval info: USED_PORT: fast_read 0 0 0 0 INPUT NODEFVAL "fast_read"
-- Retrieval info: CONNECT: @fast_read 0 0 0 0 fast_read 0 0 0 0
-- Retrieval info: USED_PORT: illegal_erase 0 0 0 0 OUTPUT NODEFVAL "illegal_erase"
-- Retrieval info: CONNECT: illegal_erase 0 0 0 0 @illegal_erase 0 0 0 0
-- Retrieval info: USED_PORT: illegal_write 0 0 0 0 OUTPUT NODEFVAL "illegal_write"
-- Retrieval info: CONNECT: illegal_write 0 0 0 0 @illegal_write 0 0 0 0
-- Retrieval info: USED_PORT: rden 0 0 0 0 INPUT NODEFVAL "rden"
-- Retrieval info: CONNECT: @rden 0 0 0 0 rden 0 0 0 0
-- Retrieval info: USED_PORT: rdid_out 0 0 8 0 OUTPUT NODEFVAL "rdid_out[7..0]"
-- Retrieval info: CONNECT: rdid_out 0 0 8 0 @rdid_out 0 0 8 0
-- Retrieval info: USED_PORT: read_address 0 0 24 0 OUTPUT NODEFVAL "read_address[23..0]"
-- Retrieval info: CONNECT: read_address 0 0 24 0 @read_address 0 0 24 0
-- Retrieval info: USED_PORT: read_rdid 0 0 0 0 INPUT NODEFVAL "read_rdid"
-- Retrieval info: CONNECT: @read_rdid 0 0 0 0 read_rdid 0 0 0 0
-- Retrieval info: USED_PORT: read_status 0 0 0 0 INPUT NODEFVAL "read_status"
-- Retrieval info: CONNECT: @read_status 0 0 0 0 read_status 0 0 0 0
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: USED_PORT: sector_erase 0 0 0 0 INPUT NODEFVAL "sector_erase"
-- Retrieval info: CONNECT: @sector_erase 0 0 0 0 sector_erase 0 0 0 0
-- Retrieval info: USED_PORT: shift_bytes 0 0 0 0 INPUT NODEFVAL "shift_bytes"
-- Retrieval info: CONNECT: @shift_bytes 0 0 0 0 shift_bytes 0 0 0 0
-- Retrieval info: USED_PORT: status_out 0 0 8 0 OUTPUT NODEFVAL "status_out[7..0]"
-- Retrieval info: CONNECT: status_out 0 0 8 0 @status_out 0 0 8 0
-- Retrieval info: USED_PORT: write 0 0 0 0 INPUT NODEFVAL "write"
-- Retrieval info: CONNECT: @write 0 0 0 0 write 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altasmi.cmp TRUE TRUE
