-- ref_pll10.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
library ref_pll10_altera_iopll_160;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ref_pll10 is
	port (
		cntsel           : in  std_logic_vector(4 downto 0) := (others => '0'); --           cntsel.cntsel
		locked           : out std_logic;                                       --           locked.export
		num_phase_shifts : in  std_logic_vector(2 downto 0) := (others => '0'); -- num_phase_shifts.num_phase_shifts
		outclk_0         : out std_logic;                                       --          outclk0.clk
		outclk_1         : out std_logic;                                       --          outclk1.clk
		outclk_2         : out std_logic;                                       --          outclk2.clk
		outclk_3         : out std_logic;                                       --          outclk3.clk
		outclk_4         : out std_logic;                                       --          outclk4.clk
		phase_done       : out std_logic;                                       --       phase_done.phase_done
		phase_en         : in  std_logic                    := '0';             --         phase_en.phase_en
		refclk           : in  std_logic                    := '0';             --           refclk.clk
		rst              : in  std_logic                    := '0';             --            reset.reset
		scanclk          : in  std_logic                    := '0';             --          scanclk.scanclk
		updn             : in  std_logic                    := '0'              --             updn.updn
	);
end entity ref_pll10;

architecture rtl of ref_pll10 is
	component ref_pll10_altera_iopll_160_d3szf3y is
		port (
			rst              : in  std_logic                    := 'X';             -- reset
			refclk           : in  std_logic                    := 'X';             -- clk
			locked           : out std_logic;                                       -- export
			scanclk          : in  std_logic                    := 'X';             -- scanclk
			phase_en         : in  std_logic                    := 'X';             -- phase_en
			updn             : in  std_logic                    := 'X';             -- updn
			cntsel           : in  std_logic_vector(4 downto 0) := (others => 'X'); -- cntsel
			phase_done       : out std_logic;                                       -- phase_done
			num_phase_shifts : in  std_logic_vector(2 downto 0) := (others => 'X'); -- num_phase_shifts
			outclk_0         : out std_logic;                                       -- clk
			outclk_1         : out std_logic;                                       -- clk
			outclk_2         : out std_logic;                                       -- clk
			outclk_3         : out std_logic;                                       -- clk
			outclk_4         : out std_logic                                        -- clk
		);
	end component ref_pll10_altera_iopll_160_d3szf3y;

	for iopll_0 : ref_pll10_altera_iopll_160_d3szf3y
		use entity ref_pll10_altera_iopll_160.ref_pll10_altera_iopll_160_d3szf3y;
begin

	iopll_0 : component ref_pll10_altera_iopll_160_d3szf3y
		port map (
			rst              => rst,              --            reset.reset
			refclk           => refclk,           --           refclk.clk
			locked           => locked,           --           locked.export
			scanclk          => scanclk,          --          scanclk.scanclk
			phase_en         => phase_en,         --         phase_en.phase_en
			updn             => updn,             --             updn.updn
			cntsel           => cntsel,           --           cntsel.cntsel
			phase_done       => phase_done,       --       phase_done.phase_done
			num_phase_shifts => num_phase_shifts, -- num_phase_shifts.num_phase_shifts
			outclk_0         => outclk_0,         --          outclk0.clk
			outclk_1         => outclk_1,         --          outclk1.clk
			outclk_2         => outclk_2,         --          outclk2.clk
			outclk_3         => outclk_3,         --          outclk3.clk
			outclk_4         => outclk_4          --          outclk4.clk
		);

end architecture rtl; -- of ref_pll10
