library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.monster_pkg.all;
use work.ramsize_pkg.c_lm32_ramsizes;

entity av_rocket_board is
end av_rocket_board;

architecture rtl of av_rocket_board is

  -- Constants and signals ...

begin

  -- Monster ...

  -- SOC ...
  
end rtl;
