// dmtd_pll10.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module dmtd_pll10 (
		output wire  locked,   //  locked.export
		output wire  outclk_0, // outclk0.clk
		input  wire  refclk,   //  refclk.clk
		input  wire  rst       //   reset.reset
	);

	dmtd_pll10_altera_iopll_181_5laf3ga iopll_0 (
		.rst      (rst),      //   reset.reset
		.refclk   (refclk),   //  refclk.clk
		.locked   (locked),   //  locked.export
		.outclk_0 (outclk_0)  // outclk0.clk
	);

endmodule
