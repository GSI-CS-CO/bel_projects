library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity chopper_counter is
	generic ( count_value : 		integer );
	port ( 
		Chopper_Counter_RD:			in std_logic;
		clk:						in std_logic;
		);
		
end chopper_counter;

architecture chopper_counter_arch of chopper_counter is





end chopper_counter_arch;