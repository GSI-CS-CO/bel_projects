// stub_pll.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module stub_pll (
		output wire  locked,   //  locked.export
		output wire  outclk_0, // outclk0.clk
		output wire  outclk_1, // outclk1.clk
		output wire  outclk_2, // outclk2.clk
		output wire  outclk_3, // outclk3.clk
		input  wire  refclk,   //  refclk.clk
		input  wire  rst       //   reset.reset
	);

	stub_pll_altera_iopll_181_arpnjwy iopll_0 (
		.rst      (rst),      //   reset.reset
		.refclk   (refclk),   //  refclk.clk
		.locked   (locked),   //  locked.export
		.outclk_0 (outclk_0), // outclk0.clk
		.outclk_1 (outclk_1), // outclk1.clk
		.outclk_2 (outclk_2), // outclk2.clk
		.outclk_3 (outclk_3)  // outclk3.clk
	);

endmodule
