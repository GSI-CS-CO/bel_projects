-- dmtd_pll10.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
library dmtd_pll10_altera_iopll_160;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity dmtd_pll10 is
	port (
		locked   : out std_logic;        --  locked.export
		outclk_0 : out std_logic;        -- outclk0.clk
		refclk   : in  std_logic := '0'; --  refclk.clk
		rst      : in  std_logic := '0'  --   reset.reset
	);
end entity dmtd_pll10;

architecture rtl of dmtd_pll10 is
	component dmtd_pll10_altera_iopll_160_fd67bvy is
		port (
			rst      : in  std_logic := 'X'; -- reset
			refclk   : in  std_logic := 'X'; -- clk
			locked   : out std_logic;        -- export
			outclk_0 : out std_logic         -- clk
		);
	end component dmtd_pll10_altera_iopll_160_fd67bvy;

	for iopll_0 : dmtd_pll10_altera_iopll_160_fd67bvy
		use entity dmtd_pll10_altera_iopll_160.dmtd_pll10_altera_iopll_160_fd67bvy;
begin

	iopll_0 : component dmtd_pll10_altera_iopll_160_fd67bvy
		port map (
			rst      => rst,      --   reset.reset
			refclk   => refclk,   --  refclk.clk
			locked   => locked,   --  locked.export
			outclk_0 => outclk_0  -- outclk0.clk
		);

end architecture rtl; -- of dmtd_pll10
