// ref_pll10.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ref_pll10 (
		input  wire [4:0] cntsel,           //           cntsel.cntsel
		output wire       locked,           //           locked.export
		input  wire [2:0] num_phase_shifts, // num_phase_shifts.num_phase_shifts
		output wire       outclk_0,         //          outclk0.clk
		output wire       outclk_1,         //          outclk1.clk
		output wire       outclk_2,         //          outclk2.clk
		output wire       outclk_3,         //          outclk3.clk
		output wire       outclk_4,         //          outclk4.clk
		output wire       phase_done,       //       phase_done.phase_done
		input  wire       phase_en,         //         phase_en.phase_en
		input  wire       refclk,           //           refclk.clk
		input  wire       rst,              //            reset.reset
		input  wire       scanclk,          //          scanclk.clk
		input  wire       updn              //             updn.updn
	);

	ref_pll10_altera_iopll_181_2yxsqnq iopll_0 (
		.rst              (rst),              //            reset.reset
		.refclk           (refclk),           //           refclk.clk
		.locked           (locked),           //           locked.export
		.scanclk          (scanclk),          //          scanclk.clk
		.phase_en         (phase_en),         //         phase_en.phase_en
		.updn             (updn),             //             updn.updn
		.cntsel           (cntsel),           //           cntsel.cntsel
		.phase_done       (phase_done),       //       phase_done.phase_done
		.num_phase_shifts (num_phase_shifts), // num_phase_shifts.num_phase_shifts
		.outclk_0         (outclk_0),         //          outclk0.clk
		.outclk_1         (outclk_1),         //          outclk1.clk
		.outclk_2         (outclk_2),         //          outclk2.clk
		.outclk_3         (outclk_3),         //          outclk3.clk
		.outclk_4         (outclk_4)          //          outclk4.clk
	);

endmodule
