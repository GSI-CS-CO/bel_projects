// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:02 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H/wd6IbjdM7tyaGeOvokFgbcMHbXW6ashVjkyufG+HVBmPG7s7WBvKqPiqQObH4t
ECx8EC/uNtN1K6a8oTooE/OKRwJaxRkPAfOZuX5v+cPXaK1Ay/dvoY0B87gYHmeb
y8P/Lj1w6D0bEqGIWLo1nY5TL8pNqELz2uzI+Qyv5BQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70656)
KXDKG90aYRKtLbYv7R+npxFsuYOYOHczK+nwbH5L1QvvrbuZpGpNSwKMxhvytSfV
+fbXjEM+tMwtgLf5kMCOuBXMysTZ220Y0rqpPfb5QZPV1SKqML5sHyGuTfD1Pqun
HMVJFejIWQM9xU9HQlcO4dr/rBUJwl+4/CnnU06HzJnSVzlm26oHIpbVc5mmUsEx
1B7Fvxi+FNcCjEOsljiaqrHd+TfeuWGx5v1EiHf3SLXWRn6tneznF20wuzAx4a8i
TJPrmZ0ZhK2uP1Pgsy7u3xmlqIkOJMIGC77Mkfq4jYSWlVYitNa74iMmRr9nWkE8
XK7maqcbUr+b1Wgv6NMKHYO7BGkPIVOQQpqOkgnXPYgfvlGdFWBIuNgHbyrE+m6n
fBFBDruqLL36/M0ZXI0tjO5Rg4TL93G32jGSLXfoi9Lm1hl7nNaFDi8K/8Sl8WKp
eK9B+Gzi/YQPDt8VMzhLL0FQYSu6EXvY0Z/2R1K2n8m7u/OvieHQgF0GJlEO0gsX
L5evOdgOMjRWqF4fSg6v2WXBLLM7nwpFV6UgteQf8yj807vYg0nTw3xCMCqbYiXD
f9Y1WA3WGWbKrhtbJwGSJ7xd6ac24zlWUG+88OTrjkjhf3YPOg+4geECUwtEAmY9
t8JBtUAPGaX6ACisHBl89Ng+FIPyjZl+foITRJdVhyfaMkjg1kPt/1oGQkbSpsaM
UJ6Q9ztTzHaPJuFdLRUT4jdTeqWVe9/RTMYntVHpazqsTsPvcF9Gop9GXimcZ8LD
evbWwIChEoieNK+xv+NxoHWQDSGMgK21r8rQu2hTCPJjuLeIe8URwbpFG2/pwetG
LJoeQ7GJR/5X2o6fOIl0Ypwqd/MDefYEzrO6rxbqaIuDV2TrGcQqMJ++XwPCPfOm
9AGkUpJVHH4wKChgndDQPHvr7gqMaaa7H3S3g0YsDaM5gq/DmlDbkzCSvNXD4XKr
OvSJ9mojxUOiWjBwakuGujMGXa171p67zYVjC8h4i8Ozexa1vCWqy/uH5EFWHHPS
DHApvUfzKr3OG9JD23CwisPkxGJXLzyYjKWtTfMgVZVuLfO9hlXo99ac44L25b3i
ATRWBjprCpDWOC6DrAqezkYSoO63FnGLHHPO4TOfC0rAZiYCYTz7RoSs2J6sFeEa
0RTfADuDZZ8FUE4lnDn64S6z2sxoOEwRGgobdskbVb0+4u0K8u6uMnbpUXkCVdU0
7RKDYv18s4bAUbDW/P5Ld7Bt85gRci4QC93FjuPAj7jyTAflmVGblHIOmPVNeX9P
ja2rNpenLvlFFMCxol+4L74te69s7RGlbS2mA8BF7WXqpd7x++zzgTJX+RcrCcsE
3EuMlVAoEy0gfAMSBx/5ZBg9nY4LhYHEDWmTfwZG843kjNwWCY0p3XqXduby0KKn
y6B3TT96I1tN5Z5xtmv1q1sfDBm2/h5Sb31a6VbzInkMI8hwMBKE1V3COGS/OhBr
GtdpcURt8ILyBc07AhiPe+ocXgsx/TA9Pz5CdJimIPVtpJJvZvhAyk5ueZ6+dft6
/kXvw4NDsuMyn9KBZK2n1N/gLi5woj9uM84+eh8fh7SMW12CNrxifuWwccxsn825
2OGIMjMPqL1O9QnnHxOhrVEbEVbYH3eQGkrpKfnYJ4dcx7TJ3ZzpphkLy9hjyzL2
ZYvXLhbWCNnFZg2B+kH3cj2JXyv41wk+Z7eBm7B4U0wjlSsLW/frkuj3cypuWI05
WYStClWuvLZcuCDdvPrRjMH78SB15uv/qD66LT+u7JfzEy6DdNQTtrZr9ZVB/K8t
DA9eONpPBU/bBOP3cd+H25xokgVGisoBQXuJpPc+Hw/t4HLeI4t2uKA3IKflog+z
0NDetE1MNQ5J6+uGFjZn0JXGBm0kD+hKjzZ3+Nz+BtwuxhTFVH2fkcFGsIx0z1Dx
NdykTC2f+lYWMgdHI7rgQJcNiDVu9GINjsHtS8aJLnJVm866XZBelWFx2VfEtyqQ
m1hKjwphxLJXm6QdIRvZwo8PjtjLas2ElNqyS9wG6e3FT0EfyvPtJ4raeBSsThJb
buFG2VXdzhcg5a9J2Zaw4BLTmwHHrWkHsMkM24JGQ/X/axJYc529I6DnrvwdbMWJ
cJYKoUuxdR21YT/cIYvzhX19wDKaLtnDpcwwD1SO+Jz3owpstRXh2I0XM3APQpEd
3tdfQrgcr3B0/qaskh1nWdK0hdKLLNJpzCD0340K39fxw1KRk0BuNYh+TzvjMZrJ
e4eLKpp1+A5LZXiInuYmDOnXihwuWU/eIOW7FPChLBIuIBMVk5pKKGh/CzfXGSaR
mCSiltvXDy9zOV2FPtszPw1PAso1vFhUiwukTv7qBrYKaqFCJzodo0hPlIfyij7X
e/QFzYUxzH52CyeIwUDd/CKbUQaGHo39gap5wniKA1uNTzg1Rqtqwl4U7PuIKVUx
LqwDLXW+62bRbyqp5ANtxgao+nL0FyOYbH9a54lPdDpjpvMD3AUCLTg/5cheS2yc
kDSsNx03MFMgnkNMyZZQwdwGsvcDrvcXkPoYXeNXTJUtYMbbFJ2dcwyy2qwhvo9w
xw1RfRF3W5L1oNKBR/omLrSRvvv3Gm1G8awH6hqSo6FiX4zE0o2P7/sxLmIGWE6b
zJ67goskEj1BuPZR+xm3nQmH4z7qU26gh4cUfWyVUMfbyNlcvOfL2BZSz4keIeP/
AZ/teYwCDAV9nUhXCfev+nmgad9+/Cqb5bhJ9kj6ks5ZqPQ/2A2HbGxKtRlHoUkh
FnQT/RSaae+/Reu2CUecd9QE/L/1eY/ohEXfQ5hZGNLSZsJXvqPjdsOBEXngCug6
NHor+K49duawKyFZz9C8L4LRlsLKSzlrS7TMdSdEoa1kuqMzsdYw5vQMAB4I7zry
UbnJiPPMxIeMU+3F8aeZs0D9fVbQaq11HdSMuBAs0ouohFKFnVW5NNSI9mEzze2b
FTmx4AgbVwdonnSDGCwaoLL9xp0JQopO6NC9ps05reZsMSnvobaIIfDq3a+r4g8Y
T/GrWNW8hAYSmG0QKSRWE+xRQbwrTKDocvXXV3S4RFRXU5e3OWrd5CFVtWYmEsvw
eK3suGJ1tXFU0EN1vtOWnNDFm2EnfUVwdkYNxa+Xfe6c6CahdfgGpJDOzU9HegaR
P9QZvEo9nkVLNIH4WqAaR9n13QqKUNn+FRM3mtM08ISt7Y4hdf66rnKnL/cuQjb5
ZIv3ZEyuKk4KiP3lDjjmsAzWXN+WBlSSdCJTI3q1nYYPyvQd6sFcfWM1IkUnqic7
LuecaXoH/anTbXze2xvUai89X83evxBnBEJmqCcbMeYkG6WxaJ/ijiNebqlUw0u5
1oL65tsqVPHt3VwvE2msvTLdhQxTXGs5Wwot/AH65LXU+W9+dEOcLDqUx4gHiRSX
IW6Fh58lMufSXunTRl3ivI9GsGbpDsbHM9QZE92RxxW1Cfp8LR5dK9HUHTF0893M
MTnVf0fTtVmV80sNWSS4r2B0hGTHZX21SXVM0Kfl5AYjfjmBek2IaVvGP6VgDJaL
l91XQIRo3fHspijIajSzs7Of/L8K6Ns+tfKyfOA/f01tueuQwXPiO42CjcFX3Mgg
/Gr0Uu7dr7YVlRdwMIflT/B3Es6QSxq9YvacQ8KsOy8iD2fohz3cMvACSDbVHK6V
WTZ8ZUNGtUUjP9cAVDsKnOuoPZ+UgheHGo3IyH8ZA6+N0uJu6emT/lBf1AI6/CM2
pgXxgpacBYNA3ZfK8S8A0177zgjnFrGAtIYQabM78vVOE0cPLK0YUCKRULrOl3Ht
ngqJUgorlSJ8ngYDdJD2geKAoYErPWxiusTdtm0NnE6kzKE9jNiaS+eUCQCRdD0U
YvMHdAnLhcUU0v76XYQlTFRQyLAuHwIhflMd39ijf3xTQamWo7glKour18YzT91o
Bj1JKRKjRy9lsTeq/b8vUnUOSmRpxTIl1s9d2wH8aqZSVFzQoR5qrx+XIEcg151h
T0haWynwpSDrwh6d5ajqNlIjIEDleVJsc+h4skbX9YtlcjOk4IypsaLGCT/Lqwxd
ofrmd9bRQBHopKGc3IfcZGR28ITLA1ZLJYtnjlpie0aEgu7UsyjX31ZGkIp/OZZk
1OE+b35673jHBur+hWEn5xgWKG8McfVFaSzGU6dxbLXjZZyXtHdzh8cg7oPXEzo9
e0jmswiE7ha9Jb3e7AnopR4UlbVZJevVFJ3jWqVT6YyN2u8/NTOlyoIePDl08Vou
Yn1MIgIrGWd5q1nqetSdBCADMDftzcac6WPzW0S5aC+lMd8aWoZnBbw4bZXe+YVT
mk9xsI55kcQ/aVxFzgPwJrkGbCL62M6/TuUbiNW2iVgK7PIIQzWm7yp0hwflO826
ae+h5IjyCyd0pmdi/bfpjj68FsQcpdoVO7S0Zbu3cmhw6f3LMOXGDpUT6z9wBHqB
n3BtfL9phEtC3xnQq/XUWomknkzdsSVXcDXLRUbHxDU/TsEFklLtQKlWswKPyXwm
L68rktAkazpwTC872IDyWlp2+yXQrzMFKsD6GPds8jmeQSoBCPF6UFIoswwPs1L7
wV7JWNMhAu6FoR96tuagefIZX8l2B6eTOShkkhbPbIryOs3fSYddDxUhgjLRybZD
NnJulQuGS59Wos91Xz2wauKgjbSauRJkeUPjdzL4dc+hfqfivGOC7KD4cdXgXQrc
mkTZgT7loMV0vtgEdoI7+VSQQRNitkC/LdH2id9HxfNvcReoKLtkqMR2yU5MZ43h
G7hdnOWLcj0AFkTYETnVxHwgUOg0taPQDQ1PjFx8QSUoebehVkVyxPY5d3n3tQ4V
+RqbiAgVAuhPZ2qQQuqYYtbB9e3gNCXAC8ZAlQBQSyIwj04KmrhyaOEogXut/y9J
2AricoVp79Lg8IsBT89+TYOoG2R60Kv5D21/Mi1T5RDfh8yDK3zYRNKp7l0qDwvt
DlFewDw2k6zY0V01+yYSam1riEIy6SC3wlVrjr3vSfC82pONLTihb3WQbAz0yuqK
thn7CFxrRCWPdIsZ9TKh9W6Wnaih1km0E3/arl2UYvFyfjYWv/PD+Ru0CH56r98q
K/IRfmpBts1lnPxqA3OmasiBLII3sLJ6qotnw16+fqT3pw7cFVabr0qt9qDRgLzA
9EJVf0t/wbKxMXPZ6hdWRzWeLcjyrEgcAgahnjuDLL37UDJvRg0pmS/gYz6d0xoJ
fYjVyovd15MDNHq5IGeACoFIA/5SV/TkWUnkgmHjUVQvdSzPN895ehYqBhJWdl1c
aNaP7XR8mvYOWtDJREGAV3rkvF/TE2BkvAuDYUnWuqBNVSa7/xgSnimW60LK1/an
i2KVjLgeJWeoXXIrgtbBxu/lAWt46BCVJtDVLzLQntfrB4Z8RplQnJR63YvssHG1
FM+q42mDZ4heRex9cx4SgduU/CUvBsptMrs89jCYBNzIVDXcSqwmjoX/1oYqgTzm
jEdjt4LvM5isZ1WoINBUnY9BZQnvtbU1Rd59BrGjD/51Y1k9H+Jn5MfKZAUYzva5
QfWkn/ChVPHNXJ3XRDahEH1y2l+zzQkIepgmssmkrei9sPYeOyGpNCOGQRwH15tF
ypM+bKGLrvRmpMQ9iBpOa77mFLu8bMUx/PHZjwbbmiE5eSACy0KaYnhVC77EUXMc
y4pZO92w5dwcayhJJuvA4KBifHKbkqFGTl/ZfJcHMiyVR9hG4iaZ6x1NjgcCeyXS
A5GIIrfIGaB1e89xMHWC+umqbWxxMS3UgEZjSBwATJ1jNwiSy+ocbdj5aodayGjU
iExXxUlj2AyPh/CL/Rr9TR2fPzbYIaCQU3dm/y44VM338aOIMmH1luEX4MI2g9NZ
mfoFBGmg/6nQXl8PgdXrW/c8G0SB418aGz5fOATYIVGwJbB4VFt9XloQNgy2cH2H
SrPZiuaN75Hj15W7PtMopphRw+BAIvnPIxoTZLvgiwcKqLlt+K1CiGr3f8OdW/IQ
IgkI8FYo3z0irTzSYDRvhQfYrU9O6PvWlElnUwbY6FJJ8Esdu6QHNLDn9+HxmXmX
+PjfG1S/e+biY9PNa/19MeQhZiGmJOK3nzjd3A07JyrofFWMJ3x6zjs09uC6Q5cS
RzdatRh4aAP5Cp+JqqWNM2j3MtKi20WET6pipG4uLQfuCaKB4oJk+CcaXwKgfmHS
nXxTKN2ymiG4B34GZ48QL2zQIF4D9HxrrDzf6IHejOCwbop9q6lbrceEE+QrM11B
kfN2rLe+9F0HZ+dZG4vN7R5LxVNrknmf89ShbwNLjt/iZNkl77OOJ2KqN/7KQRZD
zWJHhk0INtIrpAtSOxxyv8Xpwy9cRDNog5ALnzl866ZPzzB/KztziM+HU2c5tlYX
USrwQaW+2ixCpmlJwKcoOK/K24ULoBtxtbmrns1PAq+6vQrjVuyfye+zrF5DbNWS
dfxkGWXzDxhHll3T2ub3nF4mONsprNFEy8nKKjijEnvT59LHYj/wkVjbHcfwRYNg
REOdzpOxKVJTyOqAzOgRA1B0sPT90wchVWZUFT63wcZdHGHFe7w3oN6fwsZ5S6BX
yazaKK1dOx+KV7Phoq32hICjiGry0a/FGjZY6mtjgQKC5nu/6Eu9+VZu/dYkMgXG
OWr8Iya/Q5MtiAwxykS5c2ZVTLL23SVD01CsM1oEA0qxEu8EEx2ae5ZVn5GAakeR
rGrS0r22A88ir7io0enU0JR/jDpodrSsRnsqF9O/EBEAs0DnFqlFnA4IjHB6yzsz
hakzWLAAQaYuxZ1OEg1hAwFfBlXtQHezQegvKDjDMYmf0YuTbnAeg4frbBOlIZJZ
0f2mwFK7aDUmBHi71XCZ/7yn8D4swF7mZ0OWbFwU9z7jT/GOfpVFyZEDRZeDrZd4
O8IcsSZaWIXSCPonNSgcOF01ABTo6MAVznMx2lUL7UNcG+n6jsQhHm+jI2y/7Tkm
5LD7mtj5P6UsnEs7rMFpRdXwzjnXzHJ0zF0HHUu24OqMikOCveNxbP1Df1lLbB1y
OV6xCNL2d3Rsw+OpSeJSSN4Nt3WqFEoUNaYidBEJGxMCHzscDHEZyqmKea1Ex9mn
k5+ryPg8oJGs+0tz+0dzH55BkwOM+9F7xCgg12cFlwoJxp3OJeh3813dsS+11tyo
Js2cG1vOPEBwM9a3ZfUkT4t6g/2EVPph8O/Y3SakKukEEspOtQKCTZZIw9PAaKQ0
i9j92to8ToIrFZK3eShPfd+K/Sxk29m3tWORqHSOElPz7Cwf3vOnV4Cs1qe6hyks
r+PJlnM9z637QYZ6tEqI99GzMSwFxh/FPmVseOOWeAGs4qSApw06lzvVtTaZn/q4
miaK3wwqGMshK/tJkxnBWROGKWr8KlTSQvvFRjSbWvYAGayDsOKEvmoSjTu4mSod
o/r6qgpOepMU5veBhSRBFK/bPckPjEqsdbcaFT8JJrJPbd1rWt1GE2Trra0Q/WZy
k6/lLtJrr3BKlp5BdhtxaKWAy4NmtnQuLoBQeiETQIRMfyFvUfua6cntQ0L1GwGL
lZfI8NHTSfqjZWEfe/UkFJFT1/kh5eLOHQSSA/Se1+YBf8o/Gh98pQlKjFEJB7+l
Yyc92hxgZPt1e8XNf5UwTJMyB1A+VsanGDTA7c29GjIwmzLoHz2RocFsx97gDPkw
rVuDP1cILZvFIBPOOHwPqMZipQ1txrDkwxa3Kd+HjqflTi+++Q928/gsguZeavP8
FgkeReGP0WCxi7nVJHrku557pajrsyof/JyM1e04LBFsSjQ/bxiWmlykew4C17KC
GbriknV6qpaluws4JyDedTsxhmHAOEBtRhbsoMQcO4wxWiTXiQ86oHqz0INl6nFX
i6/cXttHtDHwc3dmI9oRC+BZgJJmHGmCKhNIRIo/yVKCLL8HIRyuDzADNMCIjURw
Orvmz8DVQl5dvvVhsP5SH1vdLPf8BBuxJ/LCXiqa8Tc4hBn0DJI0qj7k9pzy6FqB
jtxQEnZ++4navK9ycqNdc1keOnz640t3Y3bUv15i2uqgOqY6HddJ2SBs0/9ulQ77
EJNETEelpaiediz4mHfAVsHgRe8f4aBqEGc4OoumPmVBhLulaHW4nTllG6MZwEG8
/WsZMR9RAYXmupGbVsfjhSf6enxOjs6sqYCRKcJg+zM9lrEE49zBwnAqHR7cK5cd
h8AYV05isZmLWON/EDlGwCJ2lgV1Vo3gL+t9ixGGHwSi3TVtLksd+6EYKW15RjSz
shoQcKi54EPpn8kmxATUz671+1EYKQot5lw2hZFLMnSQzzkLyED1GsAtq0tWrlXp
R+qZcv+XgtSrlMoRMlY1FExdtdcr7he3GT3ZHA7S77MpKFWwfhpZhMycUYdBsevM
vswK78qGoJchIkRKoja+9zLaO/xaVRWn34OsrKRVjdi22gBFUZWvnyXVEEAC9Atb
sz5R3PEDtk+b41IWx1xoImYk0ZB9w7gJZsL4GnETqYPgJsWONp481b2nt2RLu9lb
vXk3utoPKA0Hj8E9AFMjjhlg1VuMIyqqgN/h2r55nzbQUZmMs65ayT/ru/QFgfdo
6E9Uz+kn0mcOSjQ3+ISgZPQLLlf4I0YRRJImzJw0Z+UJTdZf/+iebH5t1PXRQsJN
/DK6WJKE3AluhRgviJ04DDMgZ6DGp27IR9Ybt6dDbtTfKlF+e4ZrTpbzo0szlLuF
9wG7Ur+49N2lrVGIF8obtYsITrgPhyNoj7UMrnoW1ErypQ17V8XJdQmDxh65p6T/
T11a5k8pcPb4nxg1IkJ6uIEbPyEMj+c6otxpW8EyicBQAeZ4QIMnyYUcmMFZxj2d
sV/+uK87utr1rwcUupKZH087x/8tX3wAdc0nnEZCq1gZoay80WGCYvx5yav+0pEd
EIBQYVHucalLm552A3YiCWwTfAErer4wE0YESifiSemVUbmyAawaj7TxYboL8zsz
EV3ZfQX1R/wt7G7pf9pgSS8+dY2UFmc98kUp0IvYRKoy3L3WCqKw7vb61Fv27QgP
0pl/N9vdSPdQhx4dxMkoCIjyKoSVZpuS6g+asv6GOQ1oUJPvIvuLRCmjMRSxnnuz
b4ReTsHb9Kqtk81x5m78WKOVV2qRLAxzolyHpSaD/pi0206z8HUfHoeElyT46xwP
2x0d69yDFf2fuK0kCeUOsOwzcknn8l/B16y36AAqx1H+fhaYsAQ2tJbV91xbkHQG
5WtSzCSYvNvTSQBzwC/Nsgla6BOIMOGySnRVKNMeVbd5HOipNzqyd1i0+RV395ho
lOgyRWJOctYhaIw49r1NLMsy/E9UGgWwrwB2uJUldDPKz+gQkIMWcYeGuFgL8lwb
HXFrj2i5fIw40enMXXgsGUmOTwZYsiXuQe5HhP6U22toWVM31cwOGhzXOM3GjJDC
qt4bb7RkJ8x0pU0u2SSLceiOBO+x2g/lKVNFMrhBqMmf8DEjpk191FoGFpdP10cG
6QGb+pCO2VQ84iHwGj7glSlfge+1hPgfSH2MHDC1LR/qjAYKEbuuYYqOT6bFZI5B
iriiQmglnKaQC0g/nvrAh0hNFGH+dXW4ZwL00upGUTBoOeb6bWRZNBwmghzG6FES
5SOTBnHGQ8I7I2khEHl7utNoUdNzjukbv8s/Hy5JJtUqjg/+3uKv88tdHyZbKU+g
qQqeL6BXzWjSYjkIuXOswgig3/vZLgEWnZjJEp9AW9IaKImxrGb+mAor1rsHudWT
B4P4QIxeMSoQptKlE0R6N+Tv/1IuifmXAsKwrvP/3KshguNtLsPNLTDwkesNM3pd
JpbAG53protoLVeaH+D+ULJnHOaPtTaBqIrZM2akyOJr7URg9GgnEauBDjjRo94G
L8C7qGD+KdpKDeSLh2bHuyw28+vLXJ9NIzIj+9T3N/skWJ2MuDkRwiaXKNLRdf+C
9bAjIvEr04Dx0Rj9G0Gt0FfBRoUHXFZiPqg3iuhhMw0f63wMbTiQGGhQvjpHuzlg
Zyo9gfTMMkKs2WS1FV5/7lAQ9fdBg3MgUmIq5gggoHa6k1/ljEwzyMZaXY/foQjl
RMgUVy0ChvLcbcV4ZRPNEctN/Ao2ouPVmoy/90HJrBfqmyQjRi4PMrSF9irkPMJr
bxuV3FMF68UctSasEKJYiCBjF4gxm1SnItoQV5Iehr63FeXHW+gjMg+H9WfH43oG
2QRJVxYMrmX8tP38FHBYsmVSihF5ujymJsye+CBDdh8VLHjMeLeaXsRlVE6UCiU+
nEZ4ebnxWZ0/Up0OVENUVWkBqHzSUmaKv+ntS5yyMe7mcOiuNTBXGJvX5SydTJwD
v2auZlebILZXHPyGkDU1T0oCZVQ4kextbZuo1/nH22HDzpAE3fvkpFKL9YqeFPF2
ckW+QRb6uFZChWrlAMiCM35sn4+BAwpBO6P+HQVqkFzRQiz79BKk7rbq+1yHzSNr
m4DYlaDNssUulZj7hP0LmJW8JY84yIuCFa/cyeAHExvsr0YDht6v+n9wrq9VTS4Y
37RGSqsh1Drq2ybZnAjV6ZxuBWllC3X9HSiQzgBUVdpWyz12kiqjLv6FHvkYnjR9
cWotTyr77+ndvrUBlwyghhl2rWocWLoRFvBSH8jjAbDTEvCzcwstg/8M35R2pJLl
JPD5f8u7eLDEtyGFcpGRGd2W1CQaad/lREzfgqpOKVIjcYqiR3BpMJ9n2TvfYZy5
uULQb8NSHHAEkriDfsAo4zSJF9lQchEwMdIeqOQ8qsj1DY83E4Act7+w0sHZ4X8n
mI93AyYxnRnZVUhUHy13OB4Y8FePucn8ktk5V0XTOE0lDOpyDi9xRkRrHOSAQ+eN
xlKK9j1pHJh76GT/74iz96LMs3aohNDuT+A9mW4Np0FWbTlBk8BsQnHPC+13M71Z
FpD1r5CwM5WkB3KyUCGDULePB0571NIE5gO1hx5yZ6PMDbkAQ2lRemwfo3i4FVUH
JfcdJ4u/+ceQLuAI4N51ePNdAWFspjrgCIU5KlITNxdbR2xG6UKhOkIxztVFqHg+
waabV+ljLdDKi3jNK6YCHIl9eyH567FnuJC+9KQ9xQTBtsUjXUrYNT5Y2MONuXNl
YxAzmHvx4/aSuOqV6JkTQWABIegpbFBeFm8a+tRYppEdCOb9Agx198KBHR+GizJZ
d+0Z1j85ZJP4OiZC1BDfn728LghXHUkJyk07bUmExJcIvShxWahkgqGofZKb/NQa
udSKtZyuwrmlcmTAhtK4NUmltQN7RkmKBwU3ngyRLHYRKGrmzKUY4ofI75uVOaxO
GPUhj8Ocq+464p+/kOG3B6/cdqO+4vixi1qOz63i8mvY0D/ltDzCBz+szFvS89hG
cke3gILJmCo+326eglxyeGzfvZFHRS0nDP50w43XweOxXHBrLJanN+j0iGtgCge/
a7GU2hXy8MYeIa51e8fCHEoyBH5U2Vn+nP/YJpVYtW2YQuw8xnNA5mvgkHwxDn37
dJkFlAdJxSaGRlzVSso6m3PDB5KrJ78GI+jtk+1ltjV8icrL3RkcBluutATRoStI
fKJu89nU+5b+09cP3wRU/h5TXG8rCsGN3XQ0oVOaZ1MMd9A31c62iKAdEWZ/oOYW
W2Ifucpgz1vrVgc/5KZM7HGWYTAeKeYovD+zPPyWnUOOegIYUJP3WryTBj6xKbhc
FJOFJvgmsrOHd3ps8D1IolkOMwH+Yu6OlYbskI5UV9J2pZ+sWMx9YtT7gSDGqYJo
PWuZxiOEVv80F4vKRqZgLuOMS+Pw01J97X8ZE6ZatHgxOC8UdhUUbQQ5wiLVnAWh
34/fYz2Yujdgg8mGSi0kCwarSI8sCM3smmwuxAVw/I/SSHd7rpRz0gD+SI3+BBXc
LZ6V+FyiPGdwQRqtNyw1eyaFzrEFkZRvj2D62KyS4r7oc/VE7CW1RV36/nV7EQGd
anBwi+DChglVY+p5KfJvCgTOE568CB1MhV1MnG/aIJ4Dkdf3WqiRn+VJnf8r4CVy
DfGCdQtwv/hvaEFV7cNfjzHsLxohO45FFrrFz6qUaal9cNOdxthamJgpbWq6l3CS
9TcovUWUh8hXulONFiMpzmxkPOB3t6gNPErayPCXrluuBSiGkSopnXDUGOi1hldh
9Xs/xJ6pdi7ar8jBXx4Jod91yQ9rsk0QUUYWC9C+c6lXnsq/NMSR+C0oxMFM9ImW
vaK5UHcwfMPNenc4U4I1KLhISXvApsyfscJA0M738zXXWRIH+omq3POnmswM4kpt
bjNx3xeO0jfd5n7RpVfxtGGaoNDTKVemRQHgBaKn6c6e/Q2UIvsEkFuEYKmKeydC
NS8s1XBwtfg/MQMZjWslf4s8zv1BvaTbuyFhiCq5vWYfOb/xUQN7+I9Ax6thH5PJ
3Kh+hXklV2lF/sWQt6j1KMcUhZUhrsZ3s5Zuoaho9/kIihfr1dl6ySzxhGXGGvmX
tELTXzq9aqvwI4uJkNKnqNqgCunsIRQLNwl08m/OjmZSGJXctGAR0UhzU4jnX1+l
Ior8uDZy68tYzEwFwIoCIXE8lyzuQv9bkjOwrr9N5eh70i7ibBn3FrKFuzesFWbo
r+d+kxL6XLxlBJNutCWEOMhqds4YQ6fNFBf8rjtmQrjVrCc2EEzgw0DvbbqmjKkv
W1VdNdAQNvC6fjRa9GBXK9aUZyCk8hewNtB8omj3i9K1p1G8ndU98MyGmyRWz0Y5
bVpflPrn6197uYdpE68J87U7uZn5BrdHujeQSEMv/tmV0F6W3juECeiiYchLEhCI
YL+4YqibNtWX+s49jSqMg4oecIpcR1LJKwHuarW9tKj4zRt472Lmeo/xihjRDOmQ
VBaO3hkkaJG/VnQe+i1vtA+wYStN8Y39mb5Hrk6QoYYwNZ5RL7m7t8qRXrhRdX9C
iSY5sGXt0jw0KywbzBz8woXgxZ7cjaeb4P5KVDID/92CrHF7Tn461U/CEeVCuQ5G
LwjKx18/0Q8vWJxwum0b1qHLgkFmk2tENLfTNye8Aoonr1JdV8abYZx49SWT1Mtx
lx1Rh2pBNc5EMFfQnPx20fYJC17DrNBeiRiSmCof5Yrsw7zzxcTauR6zno0ej3e4
2ZJwu92eS+EPMRtyRm25uzxgL5aaebKcCLt8Q5OA7LnYm3TpoCs/F2zti+k4bFtN
/+5BG3NPFXzxy8Lzt84657A95KVy3Nl9/pO45ufGzwJBmlKuTU3uQwMvXxxD/3X/
Bvwx4VkoOtR9tABxHODmGVibc9tZIC8qXqJbqBvQPLIAOdbYiKMg3bdwH2hGJFv1
g7ltO/uXrk64cazUXeURczsMGNlfjoNEvIRe2kkIqUICDBoSQ/nMZeBToUtOk8Ep
3WQNHJR9syUbm/QhA97adtir2mlrXbZDXi5QdYK3hkdnfhcINT7z7r5HpfVp6xRf
kxjYMkuHLP/epgqbXbAOIQ8KjS6A22Ne+JGZGTajHEls8IW+bt+tUqGHO+U30cQA
9JRRGFGC+IN+BpyRG22nJN9yK/JwHpfZ5an0LeMsosQ0KaymZ8rXLfmFy8c3Q8m7
tlLFNlpOOMISfaZRTJ/Yikx4u6rYdoalUtWcPYTMqSXJCCjFsMwVrsdrhOMxbrJG
AHGfQt/xbPDLOwJ01cv+Q89qMh0fx3DZ1SKY3Oq1e7VtdCmAwAO420PIaEcppFNa
IQPbzHBY8PdeZctxeaHHZ/rBsiyWC8+R+cKqBz+RMxnA4/pM4Jh4V/KEsunQe93j
LY+RvszdAQfPabNc81HtgYgfje16j6xIlp/O2A+UGmtv/qCHBRIVBH3nixr2li1e
bAP5N+b9ZhAA5r9GVIiBIl9G6gZmOFXSP7J4L5cei/HwFTFT2i5auEB1uqYi3vcW
0X1B9lIgk35hIgg+cUM7W8vyg/nc9sBGIWBbVqLA2w0tAZ0Ksh0ZCL4VHYldILkm
aAQMYt24MyLOd5qRKYiUcZs1F7JqrhM3eOmL4okRRCLxkvVN/8iDuXqm7pxQBPwH
FkCrtrrHMc3iMLxj0H/tatpSgHvJVIzbzvV7fikN0mgSfOElAorKnAhoW4y8YSJj
uGyd4i8A69+Y8RPMCNgl637YVWe1KkoQ79L5esuoI/FbNN86UHF5YqnnSkzGQp9I
PbhuKYwA/lSC4VIZjCIEZJsXDADMn8NDL4AdLRKzte0AjXi1ILgoPAqfYxjgWB6Z
o5PwWR5ioxI9fvMgKwUDUgWfadbU53v37IKM0n45hL4O1Y3hlEv0NFbYuUXeQUtx
s16oDt5+edhNGDRKzGv/KYZbFFGig1wx4M5AoYw19ilHLEJfNFWrDGQwbF7PY0Yr
AlmEAJJ8LY6yxE35ZkawlI1rH+A1iVWbW7SgBI6nfE/KcGt6l4Gi9hw+d1+2Gtag
9iha7T+n+iUtfS9jj6bZfUGmuLfotxwA+mHGL8iwfqAAP9sRLAYg2Z3LfVy8B2Md
Zjxx9+y+Utpi0LogOlH3Te/ECib85OfzSc/x0A07PB/KBgnB6NtS3bphwKiZRruN
SnpL6caFtSsgGlIE2c3/SHagJN9MbioFj4Eq8B6AB76ZZ6rRvfnrEQ+L55CB7cCN
u9FMZyX7jBvvqHUvc27pwsMyuYFLRVIkdWxwQ2Ap6Ws4+HcPiQsHp0vm8y1lwJFn
ODL2Dqscj2oj+/G1290Q4SEFLMNNiaEVEf5ONshKTshgj4uNjBK8V+sJZzKH+gqB
nlaSCqESbk/2QvVUMI0GTt+Kg1/onyc+WOFfCN8MDD0aapnm+64bFoSBnkKOvy13
A2Y5FeawUw0ivC09mB/9z5PgKbdc2FU5vSFYF7atOibfKDv6Mm+EssM5ymSZxQTv
mfbF2mm01/RFqeYagtDsLxynzJB2B6jaV0hjmR+QONXNytTOH8nixwHEJKNeOck8
IQZf1wahsb/bjYKtH5m/IuPBGPQt0Uu0HOGpWhoMkVDi/ZyA3mWYJ5YcUeidqLjv
LZABDrCha0CZ6/tD/gsGsuEWV7jsLAU9EHHi9WinIceopcxfJ5+rj9fQS/4rPWbj
yaxw1pdVQLQHsTG+nhCGc7pLJRs0j3Kf3ia2uJfTsmQY/cW1aEPogbP/nRLPWqTR
My2Bfkwegpvf+E7zrsvIwdwNxGbPPVzEiptLA55UUsMNSmY2mM/kk6K396z28Dlc
oVUqERm1rOVhjpTcsSIVTylHTq/a77qmtUym5ls8SiWWeY8ffu4zfcn9oTHMLY+b
A/9vIRCdT7/IOKyTpozAA4M+huWlC/Cqt19pcQReHDQIpAjxxO5FjQDHee/lKezB
EotlY+w4jVz5yGqDJ4HozoAmzgWVQ/1t0fOb/eekiwofGoszBzkJugwy169OfKra
+kN0xUdJTf7vBvaa4zpy9qJri/NyOSCxoWJXOsKo6LGvSuagB0nn1P9O2z2eKvu7
XjxCUaKuxXj0fCV/LAMCOizA21uX0yuHOtGmQLA0w1/yc6daE0GGdigr09G2K6FK
O0HwFJinPEjrVuom3xReUQGxlthlyRtrbnsIgJdpMqD6aQXiKdgQNg19Zm93x3Xe
L8yoAjxEyKJFQ3souccm3ZG7rLZA3OjDTTBHp64abq5yKcbmTx/gQ+cGpFPrXO/c
GjWhU9bVJtn5QSvko81daU9Mp3bLaVGkMb7r9N0/EROXec2MpsDlgKJIRsfPIF83
ensNrJs1E5fcUFP3269JL/mSC1YoaipzrBoQmvxZ3lQ3dVgJR3GKs4I875QMjtvb
/HGru+lDvIQiyUmh00kpdQ7DdqySlVms+Q6fSoDnwHTT6afWjCyTKIY5GNpZZVRH
ndz5vOoe/qItX5KYj5GaQoT4BS727t4yk1qvSQHrRID3F5e1/HQI5RAqjEQd8Pzk
bFQxxhnoY66JXlBOg6FvZTlRIZm/lr2MV9QmzZAY3jYpyK9+WthZ3s0FNcPGoaiX
16TOHGKQQw0ztlc1U8RL2KNOavnU7igp5DgOE18i96oIlhyoPL6cB/0Fs1IndPOg
uOh2sISKCSWP7RwEZIFZB2jkt8l4b4YnoS3nVK2LjSKLsOXRP3MTheGwv1ESksi3
mNpI6aYy3BNVUNlqW5A8x1G5Y97lgAjkXmJWrtVDUIZlR5tZx0f83myrtL9fq52n
eSRmicmT5V81PpvNRq6qGwevoHthz46ThQI5YNJeyZpJOzUEC/HLGJ3sjqpvzTx0
DgoHKV8XQrHFHNnhqtwo239wrc+CmAmO0WTivQ0KtmKwZCQmr2MVodQzfI1EBdlz
qj53EzSsLtc9yv8e/HZNY9TS2KvsPwf7XAvml16JuYF8ETj3St28v8cxDP7qHb2n
Dxn5pCtGLUQ2qkKwLHLJMrcGiAZ8VSkx0GBZMsXAkdD+OuvUWKbJKEqVnyWelFFV
kI4Ch2DuZc4XVcBW8tQvTyaCpZzgf7UwPtj35H39jU4B0gAdZExKI1ltBpvIy6Rh
Y9igs05wb8m3vJQSVG6CJ3dFe0kM98Eva/N1VNjKi7UQsSgbeHPZDdoRNjmx1iLC
mXbkXBixsHz5Wh0R44TW6h/ZWaQvnLfFLnPD6gefZjTv6OuKw9htr7kxA0w+hKHr
uRb5XKeuvWnt4A6EWm8/i9NUr2ejrOM9CYKj/iGDMAkDq5cJVu2Ghhx0Qh/6vMSi
xjhOmT8cUnIvGhVnDoprJBK/2Ej4hgQKX1ZjVRFHIrkcQ0e9vMSpCajDSte4oSyu
fKp5pehZDLMnJ4q9E6kKO181yH2EnFsZHXi58VGRLSedvimrZdCzEqLUs+/lKzlD
AgX1ZCnHXKuVaQmjMwoJalkrimvr/lZ74rYdlIr1LfT+nyZQ4jbzMkHMQXXCekoc
kHkjTMHwumNQTvUKdUM6GnZ8BrHmKcxIMOjLNBrTldXdTy/06ZrA13jbWjDS0jmI
zpRX2pCRFazcnY1NI1bHw4KRbnclAFoeUg8KJbzJjmSYxOksSAfCTshtYludEIMC
5GN8Dq6+4JAW2JXj9y3gUnAkqo2+zNcSYEh2ulU+j+KmVuh/ehMMZyaNqgVEZeon
24MbVfJxluMtCIHg4jn0ONIKE1UOdeM4ewHr1V8X1BamI/w3T6gTW+Hwj6yS0iKj
99zt3sSfmNnvEwdRQJA9uuSE2DuP4JhGeALn+fHCaBBXlvvHs10l5GuYwtE9r0EY
8xkgFXgThtMpa5zmo9Atx7jDLUAJmujZwEVwUSV5ra5LKxqKFM7eeG9HkzOZ5KrI
TFZyXeTUajPfpYQnKDa4/yCcznYU7cLc8E0MIiWENDC7B6UbCme+g3GoL+C8zSxD
Y64it4nOgzpC5N+GuS3PYk5VizOJHewYr7aapA3eAneQmhTJPgWEWY8sLcMPcjck
MfNMoKuBmBmv/J9HsaowNs405agxlfKEv51HjBRUXDO6MOHbqrxm+e20vA0sZsdQ
LwSWpJ3UmnbOluY6XhMlPpqUXlFMnohzrk9HHLoe386AD+Zav/EX06brKee/a2b+
EMFCs226ea2y+8/GYDgFfXrq92hkEs3yPQqSMzImsPUXfLPHD5ss3ufXdHWF9nGM
xvWV6tuat8ABitFTxrizVWwb+WPrEaJpsFvYlT6OcVI/k0naDI5zPsyM/NXLv/hE
+sUEg+5A/aOqkyYN6FO/MewtmmDYqAFp0GgTZSOykQpFEFxx9QuP0wPbl6Blgooc
4vvQMzCRUNohtfnWPska3XYGibQr07YHvxeW7PDjBrZbsIGzJ3Ber8GBDMcxDP7a
Yqk6NMGjYOmGAnVLft1/TJX/YQzEyERMqSncsPWuFh+dxizaRObiPrA7q0YtgYrk
YIMb1w6wTRehD+ETFIHhTPOMCs5chJ3pL5DLwpJunPKq2AZNpG+/NmhpjjbVHMzd
nP2nfAOq8R7FsSB3dP5aIAY4uryII9SmuLr50xkPMnV9UYuBfMMgabVtuBYA6I61
mwblyzchLuC3im8C+CYHoD5cOheS7f9GvahWMVGsOjYhmwORywCGlN5b3fYeQtD2
0CI/1FCqlUet5wTVTnudJY4g12zYEvf3y4+jSixsxMRi1rINCyufHRv76hyUGjfz
eRBKfBKfZRiMdup1gpvZ0+mKQKaZxkVqZ5C/2p5choeb+phpcDBwPvXcROuPLMqx
9UuKOMOERsMWaO+ilzLNEY6wZzUPj/dzWg2Uaf/oWMHVj8KpUJHfgHGWvgNDUl8j
TVXxvYIa9kD++NyNGjU6xNa9zOmKxprCQ6C50RSNxK62KQ8wP7FRZRAjRDB204h1
yZAgvxrA3zvWy9V2F27lohKcyylOIMwH04qwm0jukQd9GWaBkxoMdOpk+e956BV0
gXcLTYadN8wJHoDXL4io8KVTMqX2b61FIZbkO2YzecUtDAE77TeuQ7qA6Xbsu2eF
P8KCq0PKqP7g6RY6SqM6Z1UVnN0RzyqqxsjJLSEfcsecRTGSqpUqdyzb0qCuAqaA
pqa5BJx7V1V1zynC7jKmxrE8e5kZKwqZ6SVF65LSchEv6JlkExa5jCVF/HbeYi4i
vZK5TyLJcZ+JsBMLFDIz3jrCYPvYbAN/1Vbt5j1FcTdaaXJWbsvFKd5y643JnqqS
L2uxEB5P2teMPxZLRjDJtqSFRzU620a0broGh4tjIy800yWee96B/5kednAHtpBK
EvlGUm19dUwsKPbJ1N3nTjBEcOz7odOuFWGEf4uGgAMiQpvXFULmGy7H9oa3bvBO
iDeHEg166zkgCHELnhh0/YQnydcZXURXDy5DgxA0Qn4g6/47x8scHdcgruOR5oHJ
dnpoFd508Dtckpo2mPQRJo0B+pz+ESuRSSe7E2pFS6euIWogqqHjgGhaCwAarXXP
OltBUxa19vzz+WcyW9JN4EIgQGbagDYwGmhOImlb4FDWY5pnG9Y9dP1tMBQ/Uy5z
qTR7xCTIO9G3A8KTjm7MAlSKlmjfab+OIucSE7fa8kkh7/xne4rzM8G83BDVfwGM
QD3i/A1YfD/RWTAtFoWUeopwaNS6ttbcTm2PQ2wPKGlb/NkxmfAkt93JXHPqGtlN
VC+6TN0IQtN7tycsFGBnitkPk6prjATR32iQrYuoMCsbiaLymM+A5KcVeZ9sxOyA
ahvqafYysa393UN6PHpU3U3KJlq0dlqUoQix54AKqv8gxBerJdViDFw1Ju9rFK2t
/RYcEvPZJbhSaS62+h+lPdJtEOd+2/fuM3/fi5aUusk3tV+qsdEEOhTj305+WJ5R
PIB/XdcorsOKcbeagiNs8uHyX55LuhmrwD0nP/9mZuUs2BVkc8c4OuLt6BBQ/sfc
W9OHd7fMDIl67Y5Uq9hbJ1ZjbC7ZgNcC9sLLT2OdVK1Fspb/i5kLJSV8Dq7GDFUj
w05GgZJEunu7ULiLUXcBgAc0vB704nxPFHUP52sOwqaD07/kFlozFH3O398DRdZ5
permlD5tycOuv3JuJ5TcWrfIOqzggTZeSBPwr9aZkfdh0sgwiT2ZtIZO7or0G+b9
myftiSR1KBYavc454Xpz3jilDwSzrZD5PKWr9XMzX3r1hVd5p2jF4Y9WZem5LFFh
5/v/e6iNdG+SSJir+XKgqzcvkaq1pOb9Z4pjfqnkrAwcEtgw9JN2VnnhX/LkOnJT
2TuDiCN/Xj9itsx7i+UNh3qFeSyrvL/MTLYGelaqrmuYuTmc5BZYu0WknRM+xgqK
dzMIs12XcgcnafWa1Pyhq4SyGhNG8N+uKM1XrnyRT/I2xwY55xHOhfKUq7z9XPWc
QNcu/mBc/Qv7MOK6ksqLI+JA+aaV2XR1385inZO/HDq4gaGBoaRqnX5TFC9QIBfY
WthS6Pk6O0CGAHX13kVCZLqzWVjdV50FcteDc5NUsrfDL7DgUFPFhoX0VJphWOj2
AYWgWqFyD7bmQvr+llr27JwZLnnh4YVW70Q3i9Tq2okp9SSaiEdqBwx8BmtyIA0I
HS5ltNdwV7WUqHALOvFI6Ni4PR9ys9En5eJhhVciN6NOp7yDYsJe7SNtVxgm18Tt
6E4K0dAhMy6wTJEfJH3jI61cywh8nI92AvVre13dj4yzWYtLttke2ZwH4ErhilCD
ZCxQV3oOpPQHayqxk6xettxeKAlDDtW0a2i69qb8p0wv2q5/ctKPDJg41Oq+LT/3
V+3bhxCOFaH0fEcwELEUa5sT9c1I85yyxjkxXYTYvWFPV6kI18LxvCrGX/8XXK2H
Ia2ri5ZizhgULa8/xHbzNUGZTf35rTio2cISn0Lxq6HoYsvkhvKCnTfsczbzAn4i
iSmM4s5yS4khQf3SMdIYGuYIdw39DXETWSfNJbN5e35LJ/UEiAFsAHy1KP/tzv/G
lBYG8XtCl5iGwmUBoN2tKo/XOTKUmevYyeZ3+nBmDUn5p57hKDuSX7OrVzQH4B56
IBesfJfpkLqqSjkxKjGkaCStG+cZAN0JoFW8Cu/BOZZQnRg8lzJY3X475tBIIDlE
enEo+5AcIKD6tHyV9f7z16XdpW8MrPJIcsbCKbvC1CyKH3nIkFqbsTfV3nappj+R
Z6/T3ucPNcCOzbfpKVnR2pC+JohmexDknt6zPei/6Ml7z4uFgKMFFq8hz5shraNJ
LczTCo4vMrRGkOtfPE3wN0JQjq2Rm5wlhcxur7BE9tIzySsgH4T8Lsvq4KzmJgkc
T+NaIpdVr3C5QNOx8Fg7wC7aP/b5j/Si8oeBXnZ3DIpisRBBGp26X08SyYL3/P9V
ez6FtX7dKW10ENmUQgofl6DvmUZzUKWiIZDO871+/X+olArC99Sxi9KDbZSNwhHJ
xFwNrc2vbQh0ZSMUQiTvESo/79YNjJ2QbNgELMZCdIJqOed7xpozjeqXNfbzhOcc
vu2RYReUkE44THbtkyFm+Kwqu7EZJH5hmWypSk51Suz9cU37KLbHVCtxYco5miLf
MQNF3fhNvpytTDcVO5xJ6dffwDx9prjruJaCiS9/HL7ZEdQf/5Bcht5UhyOS4OOY
jWyY+yUTl+m7Zd/7UD65pKnYAQgoK13cGBRk5H09aD34SbWME4B8oKjnLoQR81oR
ZjASSSc/mvw7j27hmCK7AnNtUVxTmY9IU7w11JbPzoz6sm1M0QvSL4fvPm+lI3aZ
o/YXCu8L0h9fN1lQuLp7MpF0EeqWCAVbgPwTck/I82gZEPoXPaFuzClB88sP2BIC
8bJmaVH0E5wH/jvUWZxkNF7Ut5iwzkmng3WiLhdVKe22RWp8ueblKJrXAVZ/vxpR
DCix691MsGeewOSuYQ/M3SCUZxhVcOO+8UPr0V5gt8yQl9KJXrfCK0ZUM8bdyZHe
774Do1bxC8sMf9AtQAbVwqP3lO3rfo7/2Bd262Udjat+ZQvZg/yFFc/T2YnwXkff
6+QzyW0i8fkaNsvkwKAley+5EeCtccjfEl/R9TIZjHGrrNPi8JOXz+E1lMbKZTfI
4Og5dQHVrk5jNvl7u+gtPpUxlti+3fODWA3q9wqCDz3mltus51p4twnQwrp00Q6T
YQ8qjKsLZqg4qHlrtk6N1AchYfjdihf+omivfcKK6tX2V4aENaNI1mUStrHi4eTT
eS074C1TuqodJfUfxoW4MZpVKgMzQPGgVfTyLzfQudwzAOBMZEIDFBHxcOLYSu2z
wQdPfbc4hx0oxBeF0PhuwGjoMIQZJQ+IBUz+/8RXy8CSodUiFY0V+QYFz9ScRxgb
PB3vuWV0C9EVEaTSHktn01WFLBYQm+adIbmCVmvR2kjfZVDBu1Ki0IrCJsTVrHgF
LvQRtrKdkswtJiQCbEAJSXt/qz2an2jcJ7muywr95zc4e8Hga3QAB2P+F7NTOaE1
kKKcpJiduHC77y+NgjgghNOZPsBQm4xGl6I4yqAXntXE3R2T5hjPP9OoVd1YHWFW
BMYJBu8MXphG2JICjwHHe5/kyj3Q1QS9ZIa7nf8129SgKFLorZgaVEO+AWBqDH1A
H9OxWX5dulHFozGWyInoODwjXdu0XBpQPrF5vA5wU1CZNsYQxj17Cg+Z4sKERRkm
LWXZ5m6Xh0FYu9ZJX+ntvjyn8ldIjg8VXsNq2W8NR7PwbKJHZfLfbRxXHuV9ZxEM
bnUf69cv82rlWlM8r/cBJNBo+fEDnrGpfeh72KSOFnY2v1RX0Oz0bZn26+E63+Ma
OULxG9ONVoP7Admz4xIIIEgZqlaYY5zs5fHs5ZWXbQ5+0SQ+EkiwyGPkfTeh03wc
pmcAKcmlkywQS+Uan68by+XPSqHt+SuDw881SevZYmSUETWDYIl3Y0RsAFVukqhB
17jYF+t8qOSEaqfFiHBXR7zfEITUmbQrevd0RDiGIgoplvYCpmTXeqaqrDnCeNVA
piNhyDXcERut/VSt8La9SiPthZOEO0kmh2dWFwkVVF3B0tYXDqYDa4lWTpzSoank
hDPsgyAkMuiQa8w1oErPs64JI9XXIKQo7qHhp9x7K8fQAdRYCyG3h5eNYUzft+wL
9jlv+rVjanWyW+vQUrpDDbk8HBUvgX4FfovmmHp0gzlVCXl+EnAa+xIFHqd9gsQo
O/Vr7LabzkkBO33nUQOYxOGSXf7Szx5Ey7fLgxGwBmjMH59DMjH2uX61c+wzddgy
Bapli95ZMm7dYU/dV1yNBCoPL5yqmFDagHAZU0uZUUlGfirPlLaD5aKjOBYZlUy9
X8EfFNJfqEz377KYbSt4qti5ygoYdBgIVrtT73v+RNke8+rwXf8D4gW9s00wjrF/
BT+hmCtV4TWjk+lMjUWLJ4NhbtsioPBVIflxf2vOAGElX0P2og1oiiEGujmlX5QN
qv/h9AzxeZluON7liHXe8Za2S6yi2afB1KP1X6DOQPoaWCt4IGrh4LRQHi7xSOwA
9UPcUPngRR9x/Pwgf0PbqjHiW7OniIPEFnp3boAyyVxwH+CUXbFcc85y+ogNln58
UitYhd+6X9VBkAYQckL2ZJDyg+lWqRQHW0MRrzUfOVi61zA8BcSHeeQ/uhnKnNFw
E+9lM0CKAe6j1HTA50Swvca4saGwbhEsvJBRCnwKpXKSq4Iln2ywKGzTxAaKrvj4
pm6y7Kfya4xoH/UAdatXX1o55lwWreZk1TGZ6jgBsDTqqFz7z0flsQJccS0f4jhn
EJ/wViwjwpZeBqSrtwO09ncG2ZUNAmFM+n3sDqFE8ZlK6fizMGfyjKherbPC50Hz
AbA96Qe0OGaEP378RtvhnJkhMnyANFc2ik7rYW4kZYfGy3Z8Mgup3iZOGvz3JwN5
bKD9UNlGD/yuXMwj1nCOyFi45v1fhM5pbpC4ntj4L66OLPMvfQ3o3kIIspsuZs7k
oX2Zq658Ubuwn9brBTcr1w7vbNyCVQZTlYl+1HEX6YijUKV/jD7llF6gHXcXDEJq
cPtXL4ce/ywshrf1vneWNNeUF+GdOY4jUb5s21j1yXEityICjc7rK/vwyVAvjzLa
8Eu7NV+Q1VoLKHocpPi06s1XOALuOXT3JAp/vy7YvZFtiHr0jnF/gfhrhWGBU+GP
fNgRtqHLMIWlT5Jtyoolj20ZM+sbyJAW6YJQIcE85TWotYeeDSLkOuZtYxXq1+y0
uuXdIWotkPmS3edBqHEVIN4jOey2aBpIJqm8WtF+7uAnOOigCkRCHlnzq5m7ZYQv
Lv/XD89y8kPSCEVrslu8kBlNh2mB50G+lvrW0Kq1TwOV8DxAkSz84dmc+tHtsJ3K
Mi9tgG/yI39B3jyKE+cJ2NCTxwHfJcdY4y8SiWLpnFwATwfLfnYNvMa+Bmq1jJV1
MC+1vRu/RbmbHyRfe3nDLXassh+RWimQaWB4xfOFPwOHCCHFug4dqR1aX0AiSzpd
J6Bgpq1dW0cMnCYcAjkrVNOCfoZbkejAKds933DBhYS41wBJyzHmaC0GqnKExIn6
C+hvklxGrmn4rOV6Zjd1yR1jl9zYvLpZHZhY7gMnKGmpTWSDD2pbFA7nliARyTA0
f28+CGmIbiX5REWBcyufLrZLttdyVuRgULSGTBrbUOzgObLad5NElsoGXkRuWlmh
mV790Oq9nwJKj/a+MuT0f6l+gqMoVv0zqaqA8ihqeBzrNj+TMr3fJAuFHWdKKPLM
Rko8PRqIDWeFoaBVqJFmWKKj06KM7kTfJb4HhSeB0+gfusoc8TcHXlElh1mS81gZ
lGGa/zTJiQMB4Igzh2OWpiAnRViwl5St8DFCTQ5uG2X3c4G00JdAMDF1mhKRodTE
dsns9GZtpCyCmnU/7uF/62/aIETbKULcUb4KQlB3o6J+RTQTxVmNvBEhKpjz6hyc
cPjVfpq7cGBdqcY4dMzCP3mn+U4oE0A623EZwpJv+G9mvD6W4OFe49fzCUEqR04I
kbiYnc5duFwmZT4G3vVBgRwDdHevL4qYYs4GvRU0Biqv7mCBTrDTq4Z6KJXlJG99
XXfzKjDNRXqIpJCtRnhcJMDfUUpTFsi7T61OlrTJi0hiTHOyipcOiElesGfwHPHt
WSsc+E/Chx3+eGFykmCC0AdFxukucxckIz9PlrJTSUhQm8O//lEfubOSWmZfXzAd
BI9aBYCC/CQy273f0qVfSSqupjEoeS8fYqj96OiI7M6hhvL7NH1dNWEWLUghmTXI
K9ghYWCe+4USb0OcZkiGttKF7oXHdHplCIag5HI1M6Mjpb/gyZ4M6cHvCgLU9mE0
fN+oJcEXr3Ur7HoJHe5LaJOvl1KZtpq8RRIbUDwO7Z9E0KDWZYTr+A0sSfFlvJAB
vGIDiOVEGhDFgNsThleh0KLrUOJ3W5+HpwCwmPHvSvRozqXsSPSXFdXHAWCJ+jIC
AMH9LwFQHQx+memd3MsJNz2lspSApg7yvXTC3Yze7zNMB1SZQKjunzKMruy+GoSP
hc39yetKBTYsdRVGTj8/kiIUiZ/mFLpAQambjTzcG2FB4E0T1xzo6vH4LxsdPXpy
iiPuuzIB7GPTcYfPAaCIAgIFGp9u01pbCoh+3JNDEJ5KQG7A+X0AQxfOox9PTvh9
/4QgYoAnZkWXQUeLbKIIGcwX2dumBGgoINO63Avwy6SHdSFzfwAqw3jAMeoHovKM
uPhfI7SBP+OU5Vtz281jDrRpm9Ok9GhFhMzLR3lN+CkSekvuNSp5+uJO3/cjstGE
R7KdA1gnKWZWR22MbdrEJLdTdPyI73op5u2RRaKWupZJRorAyPQeJmdxsnIQLjNx
pK+0unRcz/3wAjxpuFG4neiCjA0fJix/RNlzv+cWJGGUZlGFFtxiOh5kRTxlDd6f
UVtIycXL6xwHd8493cbkYIHzoSxW0k5yw8iAutj9BIdYAkGaHn1ZTP3eJuF7tW28
9vj12Pferd/LHNhV377vRbi32qWGJ0vXkUK4Ndt1VAolSCUm4yNvoX62DNwdzLid
8/M1eUr8yMzLz6Qvzy7+zZ2kf7K4MMJo4oGzddezvtKUGYd6cY+g/lN5xcdyg9Uy
2O1BHOQK00r9riPgZ+W7f3JIFlvs1+tbk3kGYYxb6pmQCpZCXOaKS02Ciemubtcj
YQI6SOXEJB1Tqq6tZH4TYQw78e8oFZR9gY15zqAdLjiiF3jfUrxOa7sBaVTNeT6V
USdsSHEyrbyCqIQ5j84QyIOB5gjaNafWHtaR9jJTgw/7VTq5hN+z3CYvn8FVcw7X
aMJtGHB6vZrKJUFsHnwsQq3YgxHhhFbr2c3qQy8Znz+5kKM1iynchTGlkYcHfeAy
sGNU2fcgeKJP+IMt1+PcjkjtwkIUPy9hSpjFxty3nXiDEV4xBkNWHAaUL4lPKco+
xawZr5vpIvOJlpMc10bIKSEhPex4fcGfddBLgQuwKsCS9Zl0HO1Gke35OIfy0FUA
mkRx/WLEG5nNbMjQOQdZq4x+6GQHsn+HyhQ6Rwj02xCSvI7sG4fOIJKXk+KQ759G
2PNYT6b+bRypBPIlBPJ8IFEQ02A9EfH9zyX7KTWXx97Jel6+iyvgi6KwYcXjFK84
xMettOiV39fvE2/Ybm4NK4A8DSOOfFpJwng6h/1OddeOqQ0OEtFG4MIgdoASytbA
YCTxEswvoMcOUfaj7Ah/h2NL3IPjRCbw3hveXTD3aHD5sHf/39tVCGIdu3FYkjkh
z7uuQe9dkVMIM4TlBAiRa0lGtjQ6zuleQA/TN8qezcnUNRfcTkTCRtCB56nn6rx3
QlMOmcy65YZds/UByymGswoPSVJd54jl5HWrMZzxkhSGRpYn45mxBPxmZUfZH3Oe
Z+6DFRxfrXfpouY/b9GX4Eq5PxugNdC2JC8+prB5If2yTGuTLxEg+wJ0jRKjxdgm
GNcxxhMZoRwYW+P7x/UYUu5CXfr1ioD2Y+RO3PemxyxgQGoQONVI6Hs2k9fyE03M
eMwKGh0BlqMP4WgSbnLTohwfQMhzH/88WZUbhoeLpY7VyDvEuSlhjxao0Niccb4E
Znf6IlnkO5eHSh12QJ4jhx3awkOg4AM2srS5WMgLRL0FjWiXZjLUxYZo3q/fIeOt
+0YSVD60LnPYdcmyqnC4KUXnmaDI1PqvaUCqfbY70jUmibwb+YcsVnWn0dpjxcPG
r1QlV7FMxwVv4Jlwb/oMPMUH9gbSw26bNWbLm10GGSn0oOuxPn+KX4NWky3rV742
en3/sP3COawcKACCm0lDKdtP4J6f/4gsg4bJqDFdCNkhKJxFZ4KJFuxvzD4MNKWf
Ukq+ahBdlYS8pgFxeUJc7HaVefl0dinac52WRLCart7bkntYJZTpzwwMp87bkHOs
rtOmE1WmQJd7RuC8PkVCjHLRhHTqfsuwAD/QZ+KR7aoBiqWFI2GfjdMYVOfdOQYO
9zK9Z+16F64Z40rwrIC/aobrqzzFFO1zh68xZrGtJIyvWhkaQqqxpBtZlWkn59LL
nbt1MvqlX8hGwsnG1z/sIRjHc3SL/JlBDTKQsWdPa92V6t+y9m4fh020M0c5wthy
853Q5wBRzaIWwfgDR4y72VsW6dRYQZnazZj0vvaDT/fiUQ+4ImQFZ9whWBqFbSdU
x/1ZLzMwMsdCCJKyFXiEkD5CzRRISUx0IQ2sEX2Z33lEHWNCYxiFAC4iQZ0UPZeU
K53byeu41e2RrrvDqaS5qK5fqb/g/5NynEXHOk9JHZX5tDZlJ73m3QjBq5wwQtoQ
hQ4aefkWYYfW0fjYP0QIAuMbKcede2omWoaw14xTRKPo27nOu0abYUg+ttEBw4N6
QPfOkW3FcLPLiz3EBE8S3riaGZQ6l89TEwuwW+FlzMppiRRdEjDlL9vAHW5ihxqX
VESqc/jhKu0sgzUGaML3eTQTKtl9gpVlr2mUMIdrAB+LEZlIGtfq2LVsz8q56qB1
bQXlbt0Aeg3dd01f7B50tWyrrARYUoW7DxV/OU3TPSO5gglD6HOMNAbEOrduyQxr
9AdjoY77JVyYsfpKQXmDgFD1XWlmX8WKzAYg9eCX+Ojnxy8xE98t0EN+dH6yKeee
VjJZt7rRi7v1d3XjAjvElp9nsrrdttWGYmZyH9hgqvHhi++0BvwOrfx2pPGsZKyb
SyxLx5xK0xEwwe5j8voRVK0eDiq+sZP2fqUXqzHJ80FGGC/eIQE+QywgwRcYQkss
YEsqPFiRvl7NFrmooipljKtC3N4OF7cSqDeH9e0hOSyCavI4uHUuh7dnjSWfsRFf
kEWgdjxXp3wzBUEit0Z6DXtccgW8NnEl6vLkfKFwpPNcbv1Hc3DeyLh7UqKon55/
T8eSW/8c5BJGHG61PJSEuLUI/Ys8QMb0AErwKrrxG9rm7uYq/AlIaPeswWk2Hw+r
NYXNTCOk67Irky1QvJnsrMW/5Q/TaXFM1AGINw5JSRYUlQuwrWumJSdeDOhUq7sU
EspcFYUVf6BZ0TuQwc6Q7IHXfsclgF8Au25PPNuJo0ZyKguB5SrKtJGLpxmbel2q
DSkUUmZsZVzPEmNvXu6OcB02J+kpw+cmYTd6rM5Es5ZVn6FKkracRUzpn/CTq3e1
L30e2dpq/uQZ0GQ+d6+fUowcLJC1LZ1qEdVXeNiKE+yebKsDA4TTsDj8yC/CR5yj
bJQW0JJJpfpjjLNsERfxjlz92CNyqOe1NjVGNygm4Zhg+D3dp29xfXpiqDO6u6JL
Qx8lNSTjiO6fLY8sa2bMlOacR53BkwmMlROFN/vdZIabPJfWyJpuFeAfkWkoi+Xr
BbQaBA4+7HiSL6C/0/qUYcM4x9HtWQ+BGjvkLPuet+7NeNyvkAZruSJlPNvi2rLy
ecVnzVm6L+g41YGTOfR2pejRa+7cSVgj7kI/E2OwX/onSGKCCJzJduJCWid/0xix
kMYZk57PF5hJooop4gjBUERv+XsaP4IJGWeWkk9nkBAKHF8NyWyqOAFPgmD38QSD
N1tGFjotgLK91wQt61l/v+RCqM+dhg38Vv16WAyISTDZetxkO/Mh07WnSxxkh6Ie
YYuwkRVT/2MLAXKt+02Xk4kYHXOY9vtIkZqA7aFvKIpRyE0deRzZsYgfINwPeQ5z
mLmsNcmkeKzQZ+vGqeCoVirKIQLSErK4QkRrKn+sIKaS7gIHoLIOyVNB6WNK14m6
/+YYIYYPnzDqNp5PD5bf37NYjOqsppFTNZ0En02RlxqVbPLvCszzA9c8y3PTooSM
R5u49ifpinhckqSTpnzeum4cB02BFdf7UfRlZhK8IjkHKAV1hoh4yyeuuMwoXeU4
zgleOSQKbbIy/7+Ckw+bRnHCui7dFRgxUjw4isle4siw9ywoWuxfxvKK5uZP35Nc
z52Wc3T/FLNaOr7PEtg1qBirHoDXOl9rfo8mlFF5sWHrzvj757ZIR0Y79v297gl4
AeZ9EgCUSZhTtX0+/Kvp2LohYwDwhc33byfk0/2BCWbVKJkYVJxZwAQ9mO5NRbQg
xcCZeLDkqvGmwWQjxu1WUCEfcwfpUm/B8GgmT+uR+qs38S87VTt45WOnsZ1C372l
reKUal/1dEYoSIQzGzF9TgWGn/tjPvazk2VH3bTCQrGuP24xnh2ayAN8JnnkKvUW
mNo73X1EClKbKHxZrsrG9dRG5xUwQ8wkSlEqgah9yP9XgUq3obj/lbV44uGfReNH
eOuEuksNg7s394FLcMFSOj6VLQoJtrez8iK6umyUsjZajgESXK3KteRLtuxb0svJ
oBGIU2hlix/BxSCMd5QMy0/UzEB/zC75nDegG9i8hAr8WKlsUU1Hj3FoisfDuqE5
Xw5StjVLLIUv3p5zIys7MB06wGpO90RpQfwNzqGl++YrPnTZH0PSaa/LMZo5N0oV
okr3MnYvbz2Kn75AZCjSrgfT+PB4Ew8a/UsT0tn5pSDPBMXgr71omYyrUL+IkGhV
d9Gv6BuCw4ajB815kDfS7j3Z+kBHN7Erb8yjvs6YuRQcv5hns8UWTNzG+nY/0ofT
NDLxtB9+CU63j8RB/j08PrvnYdI9j4fK+XxTCxRapo7fww8PJL0r3jMznAVKaDeB
elua+q/LBET2KdUS8nAGRA8Th15y+L/kC70rLxtwvozEdSCrw/UVlhGDlhPU4Bd1
2u5WvM0fiXrbdlljaUiFHfE7uJ2/XoEOYTIm58+uZ2eByFINltV4dI+AJcNLpH5V
wpYaJGrUnU5tqWxAWq2dS1lmplwURkYVBYgacMMrGGJozlN4p86Gnnui7YWsojch
e/MdvS1cY52o11dT6Oy2KZ+70h0pRpj2DRg9xK5yhHh50uDYaHncWfaoTAo0zpqU
dY0YTEd5ZdJTd82omI9wReqzFUu8at0lZrEl+toGFSRPWy+FNsw4X090+lKe/YyU
cR9efKoLSRvRJ1qA2j7s7j5UZUSOpiMBOqKNl8+k5MWLsA0k2NiBJj4xKxcEuwus
rGx8QmDLrjhLnAqcs2u3Mfn67wP+iGggGCnBvRfuXJQHktDpgtFHY5kYQ0LgVas1
BnSz5YqD71rzRFbSXAqrkvl1yoNT8HOzfHQRDhFiqmngs2DlyVaFseNpZMB+ZKUi
PDy7yWzKxEBWNyY8/YCofPZNvsPUgAtlIbU8Py5nfHQgDn2/bTtP7cR41KKf841s
cGbAa1z8Tq2EG+rwndjNxFWqIEpS1y4NejxIEjVBRaTF37nV8zRC8b8ccJageekZ
i+G6bAqBXUI/13mAESM7kNWHHZsqllire+IWgC64xnO+JBWZIxAh2WuCNQYksomr
NC37oeH0f4s5F1mwHaNC/p4iVdn84ndMQrKQolXK36jo1MceOem5NfoZ7Zb+Yj9I
UcIEjj8bZTXZVLhL2V1zsHMTjjR6wLcUtTm+e7ukOFbU+12338YPYl0mer8HfGx1
DN1eROZUXcYYl8p9LKmCiv4FLeLL4/dAkCTuPvNmZU4RXkgM9/d5reZEwHcMvh6A
QVArRMyOHxvzHZNeQUcF3W2Dg6Ex9YZx5sAJ9lMqYL3aUGcCZkJF7Hfot3nr7ouR
9VnxlEuarMx60TPPFGmrptKSboP7A7TUtAe5uG4GTI6R2V205aDa0azsCzP0ltKr
42woI/w29D/E7dT2GEMQzKaALcP/kNTPCb+7Ab1DF4FLZojsFhMbMLnDyT1J6rGc
2cb3y9FDwlqUAb68vzpeP3OmB17YBLwRE5KWrKwvsuuuL2sTAn7jluQRGaRciWPZ
0WKryUDFpZfkD+5ntN280cTU29jEs8q7K4lfN+smFmGD+KO+TGnZaHqlnzWP5ag2
AdspKQZT6+EjciEBwNRK+YScU97W7DHL6nqJJey209ArrjfiquY1mI1vZSVlHnXN
xATOL4WKnwqh5P4y3lk3hQuSA/iv+kWLQy3pDBHYwf5mODA6IFgLYR8OLuhGj161
SnJZFGwqLomMVqyx/jrO5ObQjpChytMAS2lKAIPPfKtmr8jFNI+13Edf+vyV/VIf
th/KRGgnx6tPCpIs3R8iWJ6AMU7lXfob0GCyC0MHgZSdJN9hKemphhPB8pWMr0q8
WhcZYwnqiSLpQKL1SUyd8VMbCEL2Orb5NBg0XNsADBa0r5pxiClrh38NbIUvqFyC
ulq1gSCjViPob5CcRwkammLnsdUNyvd18e11uk4jV9dA0gA2HX+tuWJLjvvXXDKh
rxeGmya0FRs7j1wfnLyRadb6dmwTlUfGftPBTVYWYjXjWjIm6AS56WON0cyvzR2C
++teFdoFCBi82u6WKCo7Flq1d+/tbIRHSUd5SDVT1SaCoTgaiDhI0XiywnRRq1vV
JX+Uazis1ax9GHlWsxsRNX88C7uCj4ZYgCX1Cp3xqdz+mZ+m0Ayq41F8np92s6A6
46/bxkoWgaQuxrXyk71h2mncc0vDZtMTV+9deELAqZNKDhxBst3/RJem3dnYYm5+
Z6Jn/IY+ESKuQl1911BFbVipsDgJgU62yVngUTGGAv1/oXWgXcgRAFxHORXFKSyy
LcL9rVLU0QJL7L5bflY6J3BLXcSECrvNzgIcpypYoaXP76CMesnvB3tQiVjfsjyh
ukkLOHrTxVhsjGfuDygmHV0UJVoNfwCfMKNZ/DtSgBVLpj9m7UwAQ4/RRLuCwm+o
tQU20hEHpuQkLvAqhkjocx7ZuQPqa+B95hYMGwbQ3OgX0w7Q1y9lV87SwCRfJa9P
1U4R4qDR/I9uV4e94uALKK5q4I3yZIFQiQ64BjjZ5HxmRBIMH080oET7s7hXtQKY
Ecpwp7vAZ2Jh7zU01Fr6ONj1riWmnifqzmjNO83nDdQZjCJ+n4R5Y/4xQoe0W6i2
r/q1qXBSYOvAgEPr41DodyoppxYDWsCkTl1Fu0rqW3Tenyu826vJEHDKHVJo79VP
YhFR8PNP7K/YUdZ3l/lbw1H1jdP0XwrWA0Oh3KAtVAvgNmF3Jh8I4RTf94CBe1W/
tjN5pLLz3vMFdLhf3gm43+t921W7YMvtCLL1U4pDJBC+EhcrX3OAwImzm052PnKL
mICiRUuPTrU8bo/zZzq1Qjde4cVxvXwGlajyogibem2R57eqoSTCV8R9HfDv+6L7
1Fgji5Oam1mxSfttNKnHweM2U08yTdfC032QjfXR4DGqtupl7B11FjAb4ZgqY9dZ
NMSTX7OZO9yQiWD5CJnzrUNE/g6+w7P0ATXt/mdddUWE33+k2XhsBw+TYGuilopN
//m+dxvu6dNojFwaa7udE60XiZN6eJ7HxcaOXMRqh3dbMtprrP8MktLVl1xTvM+C
OJ6TAwBkeoaUb5CQdjP4eG36Mu1+2uOfxCZ/mfJ0AGPDB0Z7YwMHM5wtFFNekrjZ
HsMCktDaBYa5aTxqswGTmBOhb/ycjxRa5BPfKYi7vqZakX5i/dtGXgDh5JD7cySf
mm5vDFSi9L6tkKkYli4lypkVPejP++xtjS+Q10M0/p2ZoMV404MMgXCmx8nkN500
zDcGsY3WlkT3rfE+zhr5BcdvhNAfu3aYfmVIx1hxYf6oz4PlxvxCTUj0lxE6ZbEE
MesG0kOuwD8YkFacQs7BonWGLl8zTb4wCEIZ3WOVN/l6cielOQSWzR3UwMak8V3i
UrQjv/e88ZbT7yifOQKZ4lpMwncLbrBKbqOE1W881ZXFCdFVAajd3GWD4l7m/4oP
e6ChtBv53GpZ9TqAamNym1OpseA7l8FXr1/h7+n9sgd1QCqYYKj/8X3MhKpMLHAS
UWKaKo4QCOSszM1/bUtpCg9EPqYwr8DlRJa5WAFOZQpMFA8vL+C5ExgLqq1liIEw
f+iHh4z9zLDnlmKW1Kx9gNbIwnFUgqJjvuV9dXZzhTIGseNFQWgj/lzAlgwLCzCQ
CbCO+gmmJzKwNT4N7r8HWpSJkXj/0E/FQxJfX873PbWsTFCvX+KXVRQNHfE2jFgO
f9nVu3Qh5JdoGS3nGQFsZ3QhqVoN0RYxGN2sUOjWoxGrLl1Dm3EE1P3cSN5RkLe8
DYz8IcvLneVdnfOyG08Af1xlVD++41hSzpwJbWMntHn3jw2hK2skyTwNf1cMrag6
M/AZP0RgSKu3GqNIkj8mWRHfTP/C2fcrThAwnWeCRqCsOL6okIEBkPyMKxnYOg7Z
AUMeqpag+aLkQYX73aqiaPNQlgrRgl8J0swrO9la1wEWR3QEcELTu4T4Nk0QRDOF
B6g0INRB6g8VVJSancigz7zEIbjaebcVjLBMw0BksSMlQ87AuBps8exf8+DdEQwy
/UThDeX0tbGyOVoAZo9bTA42qKg9vADFTfSkyp+yANMnJjhdBzGHZeUPjbt3RtKQ
+/Z8pp8SriIjyhuo5PVaprlMuEvTe3vOYX2JILPFWjYxge6JaVudyZnA+1SEj7x4
AFcRB2exNgxLjqGMDaKyaenPhjqGnvyiwIv5Vsfrlf6twJUSjy3PQCmbBSYzIUb0
fzmH1zlUez86qGwXETM+Mm9dnZXvUCNZqc3qWNQxFZPtPh1DPiTO+sU6ybrD6IbE
gVB+NWb7fxkenYbxih26Ccggj8l2Om9xc1pjH+WbeHjyLreXilPWh5IqPYvIJrda
HwzDGDkTLzyeQk1YipZ2UZsrAlue85cy9J9ogcJGTx0djlo5Y+CyRbC4C5TXKw0y
SaVFq6aHTIzHITZvdQaVyhmB9BHsfJFULwSvbXET36NCP6uVHfL9P9cGr6etMUYW
o6IPEbdf9dh6EUsc1yQeLrHE/TDWrTJtEjlz4drr9ZtBiijHIx8pqq3RsGeoii1H
PP4s/40v8xya06gNYU161+54O20HHgRGPFbS/fD+dxGCDUS+U2JfX0hSOsDjb3Rj
WF3zYeEFEs/u6cwfLCcHmFwY0IyoO2k3AZaBnQv9VNfhpbHfNO0WUGm6eKS1RfRR
EHm2aLoU2LJr88ioNf4yxWvjGH3VLAJ4UGXmmlXKdIkkwVGhu1gJJIZt7I182te9
2Qi1FJgsUdZB5g6z52sIW5kDmrqkoa2CsjLwq60WpOvDtXkbr/J2kCjJhOhZq9Ak
dD5He4bItayszkceBZUEifWtVR4odNwg6bF1WVFRYciGHL9gG3schNo68bj/YRdj
ZZCDhbfWk3ftEiKNDEfpf9ngJHUx4y8/+x8p99K2oiKGFmuVPGJbVdEitOi3KMSF
KJmQpj5JvKx0tHl1ZxyZCAdcOJqefxcXNzH+GCYtejQlEQRS70TR8s1/xyKA0QpT
Ou1/kVX0/l5jURCqovDH8l1Z4U4n0K8UElKs08Z/qHiynS46rnK88HL4whdmPbo/
jj4mM3oIHn2pTB5NtMOq4IC1eTq0BG2/v42d8Lw8qu6nBpruTLCff6ubhVxubebW
Jv26VUhclmGMDZ8vACJp8DqLia/zJw4pBOx3Yjf2AX0pcIpS7dMEH1f5DLc48brc
bobID3potYGYu+vA6Yn+D0hI5fl9KSKYUsduJCxkpGo+GAP5l7X5CX9bpBlnAPba
B0LKIX6CJAADA9OTeQaAQTKc3uGXL7rc3SQo69DyhAngAPZqQyD8sx/nyzzWeBN4
pBggWUDhrsDMBJZmTU0E9hyM+thVZku+G+Xu2UK5qCS6p04HynAZPbcKXdgJhBMF
US1KGnh+Vq3TrDWQCSc7Z91pEQ5l5mkuVPvBeZwoS+ss98GDhVs1tVFabunFRDGT
GnKtBFdPqQW3RoYeVZrDBJfHd3pQ8NUjOJ4nDJknkfdbrg64/RMH1EZusiRNkDVS
IoMpeatMGUnzSnLKzT5FTcj/IWYdkypZCPfRNMCfEzxiZ7lO03jP+yh0X5GJiCq/
7LehCbaBOEsP3i0iklZVZLKwpaB/C/nrSSoTZrwh0s/L7IUfCWCY9GMDlw3dE992
knqJs0CAGkzKippSuNalN7tbZvGd+eKjV1F8pficO60Y2fiY7bibhS7UB7gajZ22
j1gt6OIIA3zKz4daBqAhBMuSrYy2VXbY2wFDR0uYZkk+mDbZrhyV+aMu23lAbtJb
Dg93wmoywuuw7oJixi76kRe2CT8GC4grWenE5pfO4NhH2ORP86Hc4T1jINa9UnCH
kc0XpxvxJJKpokpvFO+oNmNdbqThI7Lcrlc3aUoYS7HF4mFziuXhXEsjXQ402Lp0
R4tC6lM/v/WUb/+G4GXgBihstlr2LB4Aj5LcAW2/ikfmtj/2NNuEX373etZSLhau
9SLUztDeC5GW/Kc+aB9KB4eSKy4pdyQPiC78kFHL/UL//MIs5+DVZeaoAG/WBgjV
gAix0XnlP9lNwy/NknNnO/v6fiC+1l1y19mWZOZU/euq0gjJSwRK7tbQ9g1v1659
QDCbbccnV5t2XUXi6Pc76fL5Gdwk5s4nPNFyjKmHZexDTcwH5y/Npsf4Xbw53MkB
/A+QqU/+U8FbWPILJGEoCpcsJ4hVr156BpO2ux2QLuIm+9Eqtw4vKnb62N9nasmV
tl1FrNt7HpnVbo0/M1JCl8UdfCjfyAw91yj8M/uo4ce7/9SCioZqZ3R6bp9F+m1j
Ty8BSrDz2at8oqM03Dasl/OCF2OY8o/QClUiLRwqEvcpgSmlMB9632D7ZQTv1QSr
mgCToKGpKIUCk+fB0ZXe/cy6SDKeIrJ2kqUAj6b5it5Gk6meEsFBNwsvi0lsRF6g
SLt3Src2WzkTO1Q2AwOHdbAtfolS4iSOo5ssyutrJVlOUCLm+O9TWptC1D/wAlvw
sQFU8ZR/T7Ri6yAIO6IEYWJ9k6S1Ed9H/UYWnXnSzv4lI8sVRzzp/b0zIB0Xq5g/
Rd4VLt+Tl9T12SKp1VoVKufnSIIZAThnn8Mgq28EPH7f2tmLzusKKqoRXECqBQr0
/PPdiTUUJs2Qra+MzPW6b2w12xJ3DED0py54A7rdg0Fgih6xuVzWNWhzqZYQiPUH
aymz0rCH5ie9ogG5DQVDrp2J+BDPi9E+nzYWw+FEDdB5wfG8kOcXNuvI64B2Clho
QCMl4tt0tWDPiljUxGUfePdiigo5T5oNIipkbUXZ/myV+QYUQDdos4eLR+ABMDyL
iZpJ+CTLJBUHaHHh+ew8p2YuDwpF3dPXafW5ZDcOs66nCHMuc5beLsOqY7uIgRVJ
9NlzloXi6IIoELH3p7EkL0RNrgihbRhBrSbfr7awjyYzFAKB7ug5PJvdyyp0MXu4
sUdptkctBz6wH6gI3PZKhELAp/S7CWnHvX/9C5OZJf/gGohyaDDorXWzOUpDlPvw
PQZqsNMjX/+NjU365n2qLfLFvSMcBaWU+SVyCTE+7oIPgz9YFEfTb5jtUUrFJUrm
bB/B3L5jVx4lmzHL/F9Y3yc26oYYVOk2WJ9a+ASPSG20w8eBcGy2MhD12gavGuem
gN/br0JSzP8mlGC/WrPpevXbC08SEQ52/tnyb7ta5GdJLu+zJHUzHnQBvhXjDKtQ
1OiCwrgKB+9JqGiaUF7CKLhAXwyJco9GCbLjWRKVWqqmfUFWRZpuZnkkvgme3xhO
AgjaHYDXoF1adJ07dQVDLfQYYAnNkBNLm7PBcY8ut07vzjF1wLZWG0kctOxeiYkd
EiM+vcnpN4IAtsCy9EvximqLe5aKBDHAikeEsyfFKYNrbD5CDoeZreNgI22FTE9k
03l3hyz4fl32i1U+84QQry9ePgghE4achsBJcnX5kKDs72Xrqf2CKncQSB9j2oAH
F4rLf8DgRda2v0oIfkzNX+GFONbaIea0I910u92DeVuz/x73RAHx2vIcz5D6QPV4
Msj9dCJiYy5LhGHvoW+9pc4jka7s6BfFoE1TCrgPRqTtcEdySa1zQxcb6kqVHPq+
lkJj0+t3JjzQ6kl/x7hkjpJsuth2xpb8OSAFyWdUAmdsiT/zZs3zxWn4wea7Ab71
dEkQN0XPgJITGM9NdjwHFW1MRFVALGGREcuFF6BQuD/TOhbob0ZnFowt+EZvSOhc
ATh22KaoTsUY6GUBlcvwbR04RvJdgNTPt4LivTM06z1Los0uFA3fQ2vh1WVA17vx
cN3+sKnndXSb/VnuQHgeuFq69KhcTm+4evSyT3bYQlho4LnKIU22G+08E2ANBuW7
HqadfIwCV9aG8l9L26rtCBv3CMifpHtMcPY9OxVY7wf3kd/VUzoikGTwXrPb1rSh
HngRGvctbiGUUlZiySrYoRCXaFcoDCbzY1TyCBWxhBz+wnmWTcwFscpjcR/qBmhN
ZZr/994h01ud1xu3RD+zmCiAgf4LEkSBzJE1K/WWnL36/Pu05CGl1lWA61UpVA4D
MYd3N5zIg40Bh+iQG5jtPt7p5HPHawd0l3j0qmnufmkxwOLNjF6s8caKuL0hNUCg
fZoLnSQAr7SPTNDOg3Mr9G88l9CtfoNuyiPo1SmSLs/f6kWjUsQ4M5UIx4o3w0pl
OZjxwQmeku2kr7B7DTYG6ELMWSSaFpRyGi71YXeO4t6vw31bDCI3V9WjQB9yr9N2
dbqxqT1bU6hzGGnEMMIuPvFC1PFXr+0tOryH7Rfe7+KeH8wERKaVlBWQ0lfCgccG
TZRtcJ7exg5/XZ2gVSUq/O3PWfez+pmxEPXUzYeH2xS5zqjuMxu2EtUmbThPQiEc
HekPYO7WUbSOoWBSN+TnuOLe99FvKKF8QH8O3MxASaGp9WsTky/FqK6O6DaAIhbL
iYcIbO3Q+PAPqaqqKw8D48UOA0ETlygXAz7b9nIqcKoSp/ZVE2Bn6Yc+sr10vJ9P
RSykufR3ZdRcpMjb90wJtzCKVoLXsLcn2l9uRL/PFhvBDv0xw8CyjW97GgEtmhI4
JiQVLKIxbDL+YNIojqCzziJcUHOJqfKSWsMh5VDsHU/oMA3Z5Ioq7cFZ4CLy6x9K
eb9LyGNqOFWpU/3FTLXF8ZU+OpuYUj89c5lfsBinjFWKlRTbSpY5iwKGthYVL4hE
57qTR2Z237gvc7mjp7nWeCebbZaDWgo4G8+oGQ7pUzbDwr+tYidQxyDdh5clXih9
yNP7k0GJsclZvKfYRKmV/7+EJB9Of61ikFD3x8djwkEQTbTWL6CJXQm4zXe2Aomg
XWYGoVXjhbUcWxbOYhtKSkK4M24e3kopRcXzUBxhy7JkeAP1yglVfuituWTYixyv
l84Tpv80jFjZuJ2943KELNY8xACFAOBsltdBvs5oT83XYbuYHvp09sqwbBoRWNtQ
QFmUZjGLMK1CXupz8WgEHzRIrHIYBPgNSy+A89x7E9k1/S7M2IyB/ejdYfw57t2S
w2usT0Tf7PsILubgymAMqBP7sbMmCVGn/SzZpEVRE1kj7Km20Bw3lWVejolFDZHH
UnQDy9RJX+tSjJEL3Mg6S9dJ3AEzQr3Rgdp6ocaDgAKKdlVCYaGzK9W81hcLxORz
JB27vicyP64LmMd8M2ya22FpwEfAxXJud6ajvAP+yv+PZNfBmFvo1edzm/VWOHXk
kzUa8NGcrqqdDvcshEICFYquSS4/q1Ze8MqQdoYosHJ92kZiYGYs8qY/ZGozXLYd
mB98WRTyl3IeUSxnLg6X12d676NH9FrHixIH9qR0SxsEGcmXZLH0RUPx+Q471UsD
zjOhH0jzWGaZthrcfmf35G/g8fdL6XVSJJ5ktqZLgbjWud9q8YVk/pzCnoAFCofK
gBfyt+9IoTkGywhjcp0FCQxdkb3A/f7CaxMBbp6HoRrN5QaWfq7ku3OzAAVLZRuo
rL0l5lxko0ZFN9E4wrOl3MaPE5t80c4M+kc91o/pDUDZf+gWI1GIQOQ92PaLmYDk
qLKHZ9Fu7FffI3JSHELfAimYFkrn9LMb/euQnqMXMl8jVhrOXC/mClmkt3JVj7Ur
yz7u0lOuTxg3gxoNsGBsBpc8CZXL88BM2jT+Z9u38vHIUOnxTxGgHceEwXvJID05
VkvwLYQSdVkA51sIvoFFbuzf+FmebF+n1lBnfmEaCvUq0LPCET9RT3wraTmlDmnS
1rh3kHk7CxUUc3CJxj0hmZgqWgqlwxpTXytqkXwA2+3Osd1M2X2mtVyXNguHwtiu
pND8hUr9Tc6BbkY/0SK5fQbfKGptKO/42c+3Pk7KnJ4Uap9jCG1sp3YyA51BHqI4
aCCzP2D/wUnXA0hcoGYcsXY03EImkGNi0+zC9XaXKKXNA1kf5U3MtNJnaUFY8xmd
iVC+HfJZ+5nBbn7rhvj4hDAbvss4MNK02gDWw19ifwUkyz8h+v98ifGktl7BRAWM
DmeQxIR5NkoQ5taTYc61e80e+B0fXitLEfo+UR3yNX0GeU/pxLeR4kwfPawfSaGo
NGweoP7VDIhzRxWhtX8SAxyCdw7Lzth8/LlGfq6zpT314LvmM9+u6tT0xsB3iqcZ
E+D6co1mygpmon0GDErxMhUfvT1rbCktnOA+P/aXTNP9D3k+UJ06OnDSohiXpTBl
69DgNSzSDE6+90T1dHEk+n+qViZOQs27Ld/MtM6mFIHOynU72PIXPtVcDZUeMqdm
WFN/lwl4JA25cczmjwJLXHqF8YHiYDdTXS4edTNHarWUxguCQ4L59gwBmE1/SC+d
Blh1WHAdBNA50pA2R9cOLT9n2mvThWHiHtaZw7Pyzdf4dk+5Kf0VbK8j9ZONV8SL
ZefUOSk0BjFT4caLokycvNvpUJ1QmZ0HuFgib+58boJWNV0yARNtrp6J4RIWPOc3
rOAPxMhYWkrGPaoIHd2VBm6p19yCk2VnGWXEwDHhUmWaKN0anceWYAlLyK9YNU08
6yFHsvIbKEIeAN8qUisReOStSyRHky4+PXuy0enz5zDMTJ08pMu7J2xuVylI3QXb
zO/eczBUNvbULDxfAdtYjbKEjXC7ztxuf8mVudaF3GA3jJJHeDnfkEgfKFYCi8/Z
2vcyuBril0aqNBjTLKKVQKgEN856X+Z3D5KnVu2zjZm3H/bYUXRMz8SXce5lYW9H
13Mbtpq96aPgZTv93FU/fyn0H6HYG1De2ACMigxmQZXwQEeE3FCAEec22g6Rf6vI
rQ1ri0MNisDfagnUVIcdDiflD2DLMN9ZdgVWmqyGQinC5MCW5/gqQbz/1Kcw9nyj
SB8Q7ThT1eMATLDNl3h1jnUe8j+jaLTdW1ddPWWKH++LVbI9rdNXRUiEImCXaHgh
scHe2h0GHew2p10vkxXuEhvu+z5NkbeqX213bksLeCYCFi2Ojg3hOaVVe5E0sxCo
wqrQUz/mNsI+YZt5EWjQDVnsSkDKcxlAhswfhJiyFVZ7gXCGrR+CXQYTg4vDTgJ1
UVFVp+ir4fMhrfOEtRZ/n6IEnPxbv5KdZWDLhnZUQpwDPxXpxI/q43LtOGEsZ7AQ
bKz69G3pAtgjTiQVqI4NqkwbLboAfX10j5Z/eB4vB5PGE3TosrF3/mCiQqJRFA+4
PT4Y0wZ9hc1ZoED/EdmqHRLfpYHgvMR/WvOXnPI0a7nMxr76VxbU97ss9k2sbYKh
BPxPihuQj9pcle4wOQotmeqJL0pmfFp9HaZknGVAq+geuN+iaKoLIFW1c7YMN9Fa
eLQD60H+YZm6xgpJsKLMEgkf53cG0Zqm189R2GizAhEA9quzu9h/c32hBY/VyqT8
V/UnFUqVV12uuKBXoJuSGUnKtXoiAwgXDFXcg7NUnOuB3xnzXiWkGHzSElTvgzBZ
Rp71Fc9g6QA0kB5Zv/7Y7xzLhuf/07F1VwHl4mVT+slm77MMBKIczOLrtKZNcxdF
DHos5047O9QtkDhfYXt0Zi4FnYN+cCOfHkPHelox4sP1TmLj33ChBA9jAgCrDkTe
hgNeJ5dgw9w8pi9ggDcRieLG4YMcvWuwIO/hZ2U47qfUjqX0wknTMOHro1PjsZ2y
LIDt9OFGX3+kiwIF6ayCQmXZcWzLdLAhVXWn8IY43BXRqDwooaHN7QaIfTtiI+bV
S6OQiZjYHclQZAlgWW6onuRvjziFNvVMbStlT708C22dKDmmrvIDA+d/etNDPj10
63Z0f0j7CTqmfUaQgUhRR8/QY9fw/H8tLsDe8at9ruxuIwsCUV8PjaxR/bU4jvHj
g6Qd4OejIyBjdI6F3D+91PUhKLwKhs0VtQlp0Lm7E+oZYSMo08hOdIppk9+a6/95
ZdhX4z/EtEpqHgKIYxBIy0mejmhIjPzr1X3AgLcJPgR1Ay9GMU8R5KXKv428W2kM
kBsDzJFX5+8teEGbXkNztcRAp1QqZESYHIgE9PEk82oe+KfPLwWzPOPtKSQOq5ug
nt6aGmEYmWW4+K5DmzuKnFERCxZc/Vb6McpSTRKFLtNf9ca4ivfYKK8U3pJUwcyj
TtPMa8lWmiut622AqeP5T52A2ogz2l4MKBJUnn0ldzpvzWYIS7Vs4tCYpOll6cCW
/yE/Dc11QBDzAqjXNsadXbpBHbu5iQDE3hc3wTcfs8IMIZtXtq8HpAY5YJzMZD5z
bydAmGsiZ8pdOLaPLl1JlIUCOCDdYZQS+G3C2kQ+kKR0gq+b9OGu8vgONGweuhw8
++vDdhJ9JexXS9lxJDXYguHN8odya6I91l5IBFeW8IwBc5igWM3srf8wViH3allN
Z2e1+Z55ZuVVoxXt8/0fyZ07J6TFmq+TKuxx+MwC2PwnL+QUKSS268MV2fZdzXWA
OUoG0XgcWYRddkLQFh5TQVyTCoNtxaJxtX1YaXw1noIX3LwuFqWyTHPO2pS3WV5J
mdS3K/MWIojYIev/vS2bNqgbpQExPCElq1fSds6tOWqlwmmRBQJVLXM3WMuZYyKZ
e95sPMiCraiEI6Fv/JURYVAuWIJEhtLNv66e1f7TbRqNvgfLI+8zGnNCsDyGWQba
WtPaUk6GhZ8k871d7xnCe/+qqaEH38COaxThfG9cBtN+OwBz92l3fVrHSpGAbUWL
jfzVriiU9sjCrbE3ex2vx2s215MNjDnD9AEytjKAQAOsyxRiyjMb+4+Kg1VTKhAr
ntrXR1aQgNcAJaclSiQLxyxLkp8rAQUsHwnnFWb/ITF4MsfxocWc88nLpcXFcea7
VdKTyHqG6VX4AoXMFsUvIxZjF3oXeUBhHcZmMPPFXyDw6RSMGAwjZ/DRdsGEMhX4
MPwVQxEe1ww0ltlDKYjVjeO/8ixkI/G6RLQyaF3pKTgI5jc7xs+LrMaYveuZVNlI
RE4pyzqfx6XrrZaFWilpFtpSGcMOJQKOQv1Sk+ddSKJ4ZLnvKzHbPs4KwfAlGE1i
Gqe5KeDxAEulGN+jThBLhmN3J2c10UAI2ge860ONCbENLZtvbaKCD6j3wTeEBiWL
oQj+A+zG1UyIiDuP/2FhU22y2JHrpIGTj0XJSUo9A/6EJZwBzvXiBovU+Pq7A0Kz
w3IN8e/1zn+gfvXuuljLKG59rSmBh3rriM1EVEbAhoE1FAESgn3BTeFyYP4fgROu
7q9/n12DIwiGL7IFx2rh3Ukbif8PqnrusdPf4fVFas637O4LvZS4R0MsHGTE8n0i
HmJxgP9DVfxJNNWMYIkVATo41Ol2CWKmqA+1+tQjSLtGTVZt619HKCk6rCJU5TGG
e568lxu82WMktOuvvAMrBl6bEtfLs0JuhzwRUPKkqdvyFbQFI8pBWvqEcn0eXwuE
6/5BY9ebKCx2iPV4p0X5aPiW4AbHgHocPP9xJHszxxbPQIpccRHQdytWp1+HQ0wz
DGJfecGkTdaDzIcu7KnLS1FmmIIrHY0Y52wq6j5hI5KmsHUtDqR2Z3Afr4r18aiJ
qEi4TWoB2GXpIXB/hoHPpOIN1o6eN7ivTsu/tVbFAkQAUck3sBmAyAupmqI5fvic
2D6OvjQAtI7ugASdNCm8/1Ifi+WfkHz7HMumIT/ho6hb/1r6zE50+sN67Pw1hTo9
1mXGCKSWA0PkC0VKV0DihS+tfCzyZ2ndDiotygZ7GxIzlo3jOqK6Kbd8C+dcUknk
vfV62WCyhj7G4kj3T8GIBh0oipi1YGbL+zV5VYAQVxxo71dMWq5DungOT5I5QjwN
D1zDYZgxEcYqITk17xUQbgfm06cMJqVn4LUQxmCRpHkMGlIXqS7ICZ5QTaDVk+gO
LiD+/sWrWO6wquMsgiXLz/FwiRolXphTVsvAott87HGKIV6b2tVoYaI/Ez/b4EVG
CXSW9fDFan5AgF5xA557zkTvmiic/Fy3toiUcFPfKtAm//OiF9bmsf54fG9Zh8Wz
rKwWabeXmVmFI3kbW+8Ow+Gks1kNTuEqeFZUrOayOkOZBU/hN8etjCfEX1YCs/NW
YnI3M5QLgSR4eNNO9g3frvmwaid+6/71Ztnq5vdisypUlEGU+1UwGuOP9z7oJ1v+
mak7Qmk2BKzY07xtjw/oFq/mjgfMocy0s0ueSqkhZjbBbAxLA+8Uq4wJBKcBm+Hg
CZ7zMYmgNlosC4Myf4Vptqvt3Zn/UtEgpCC3EQVPhh0/ffJXmqEtA4XjsDCGAt+7
R3//nI8vdG8MJtfo0Nj0LCY/0lvf5aSB94X4wDnwDX8xWvwUwGZ1xQmkcQkDz6ji
dE9UIq75EKfEmwMufHG6+RCjLVNG1jwrXngkO4Qk75RcC/7dEzy+kjd3ztfC7m1A
zAaIULHwYtGgwC2mgpZEygS8JWT1U1aCSdDHeoveXHOvl2lGpgOzGSCfSk3xmRe4
/DwHIRceM6CRgqva+hp0XuzUKrMsx0wma8luMOQcMR+j3YuaRfZjNau+Id3rSOdZ
xqWvea4nPPgnJUaycB5z45huxf9VOM9XKlE419AMBY6mmWLagpUSkzsRvBu7BBUO
MUi81mwEgPcCWCpd8bBfRvin5b9xJTEvw3XkRYoTmhGSS0lU0T2R6GiGwPrbDipt
CgtW0mrTgNQZhmYeM9ioyzp15dViUfDzFUbTJLLYaOQ+04I2ylS2edNFhHoTz1tO
N5wQc5ZoSPhLtqANEigoQPGiceIk2Y+wEUksA4G5MhHQcHOYqpcrOHXti9XTwpjz
xmBjRTSv5glv90qIvEKSURNR7/Hq8KCUXKlcQXxQmTrx2WKfEQ8VLKjyok/VhE2J
1EObwBQE800mUBg18FwFqJSqYZrnXNvdLru311jn0CZ3Yku8YIc52qw98ir7BGNB
iwtUDADTqZXXD1KXGrRRSsp0sT1nAxYmOYi6aI0+YGHpKUrIqYg3WHqMyTdHcEJA
B1IuzuA2Q8HCRmvu9fUN8HlDQuzYl4jNmTyBSfBD0YkBApZOOLZNpCkFJ6zMSf9p
7yoZiNt9fimOHCMQL5F4pX9TxATmM300oFia2yvDyqtTfXBSppHUxfBGncGUL+R/
7KakbVXjVcB4JyjeSRhv5NA3NqiRo2t3BAMfDSlkxJSoZnS/9zy3lY3/4jwVf8yo
o82GZYgdivI/AMg+2GMDwO84tLZgN0lnG7ZnsF++uxWBgmg4zsQHc3ft9KY5ZHIk
QgyED5kOxsiiVFX+1fdnRv7nbPZtz7lOQ1x6iJriukaNwqdzWzfxT0ZP4JgzIezO
+ed2giQiLUSwZyCq83xQE+qlZr+UNI6EQwA7T8iqMZkxDDsn90+FKu4CzIAK3Rok
dCGdtlAJM1vXVvpApLP42fLMNE4A+zhvqhAJtCG5nMZA/BOM/CmU+qap8ZVqWcuH
XXpABLHDtK+dKs5fah5zy6vEMx+IaBxG6tEjI1zbLLU+eHzztbJIaDEkvKf7DrF5
d6fvMCdnNmd9EMrcipc97dKXc0nTPeyPoaY2x6flD2Dtlvj/MrHLgAYz/sUcRfg5
U6skxehucrBmfzAb+U7g0uPDZl73ndkEHp8IYhTOr9y1B10ApaFQ+4z7ysHGwm2w
1dRe4pqBg2XjJUNz3dBOPpjzBd3/pFUDkAm2d8jFE3JrHEE1xIV3zFd1agIaCwhO
RgBtqb7SvZVr6UsJTkUdCqoZ/rbarA1fcM6v/CH2SHs1ENn5+9rb2hQXrbDIHBRq
MWhqECE8dn+SopNFWDxfrCbFTEfzM9HlB2kQNWU+Zpd5PL70VD42FVDCn54I6iaF
mdbSnraWlMexD0EWLPgoF9RiHhHgFVqSMuBJGwIoqqZ/B1gsUje1aiG3qN5LcL3X
FH2OZHvQ9C5bLtFQSc/bP1MgZDUeznhMB11we6W2M7epBF6+ZEiZ9cfkhDwimEss
1+v7xJkVip9ICsNC+AxfVNTHrIb5CROOnjFoZjX+O25uHMQHWewjokbnW/9uEAqt
YqtBJkCqcrMsrEPmmhXWI8eioKMIRZ3wNN243wuU7hKItiRkKex7BLUp4DbFGIQV
kluxvKcAT4uQ3b2OcXZTiRpsQld+EniuUzYHEXCdgPM6yaqmrWpOVOxLmlP+6lW2
2lvBijYoWcyDZjJQDhfwbYdOXdxCZ1Mx2cV5tgdSBDHBr07Y8bOX4EsdSWY/uOqD
9nHfvndOlSNMVu2RlC3xqx66J2Ye8huwPV8Q+WZzzJdl1a74xKGD6uukPBwI2s1o
sUe1TSSx3BP4LO+oKI/9QsPfHLwQ+ZInagfUhTYclwg0/2LvljZy1SSm2T5KUbBi
CJYOWprTfh9xn1lfDIUh6FkmXBWK9RaNLuF2MKRr4GIQMicr4d0CnGAgxyyYXkpQ
PhSn40GkNGxl0UH3qP3G/N8l+FS3o9U2gW0GfWjetId4rzEdTjpk1dmPTAbHxJqo
l6Jlt7yAXYyw5o1WpW+Bs5zsGnQd1dzcYS68De+ktwKYKKWBO+G9FGj108oU6hs2
JrDWVW4IlvgUaQLvp+y+pO71lzRVXUHgFggyXgL4igoCxpdlz2nGIEKfBWyYRC/p
5GO7Zslgw29yumsOHoJqqfK4S99CpgY8Per4opb/fMfSxzCypxTD0oh5pqRFW7Np
KKYdCqmBLw8oqg6oYx8n48YKbqtOjZrsCs9pnXmR6opxMrpTlVrs2EwVtYnDHB22
YBfhGEhJ97HH4Pimsw/zqvP2qPRc74PmkrWw3zqiiKY2yR4eGEF30Ujt62GyeBk8
WOo5dZAqZUl6S3HLX62LBBnphgSjCDVR0KoXt08XN73QzOWrK/9xD39GCJ/spui9
9weHugjt1VACwbVsAVb9zYkbu+A7Ntlxyn7Xgz0nUUerJ3Q4iENAhL0a3Vt6qsMj
DyyYS66pUDXWGC4z5EScLrOIYX8ZRscFN1eKDykO6XZp3n6x4xDbXEvfmshyuZYH
k0tVI5WUg6w/riWQZQw45YpaNlDxNWfMr2V5c8gZbItLXpexZJwbaEkknFvoBJDR
xbW11qQVS2bMUH7F5U4SRDtdazDcvd+hktyPeb+FRWAM1oRv9MCPvwruk1vdISE3
k02fUJpl2ELSTNPzcGqG9kmKwgIZur52uuFR2JDJhAlWkUX+uf+hA82/lsAotqvS
LI3ZR9C+lw1bcPcDdlW+qKtoUnpk6dVTtLHP0g/HoJElAsdoQ6rJ6ZhRFNoi/0CR
FOqUoqXKiBm4U3UF6WoznQHdMz2f24XEdN32hHefo2tCrSwgy+otwvbYNZHm9MWT
Xi3gIpiAs7cL0AJ/sTF5gmlpeoi81v+0sVmwkB1hlIQ7D9O7RY5oRJlUPx7QTd9E
ne6QE05ayhFLCr9AqHj/LOrLyl2vt2CTN9dKu3HYXWrYnxr3ce6uvUhcDwtZQi/j
OvqNM/V0j86ZVEER3jWPeTtKdUe1GSPm/5JUY3ZnSP8U5KccAT4tTRRMj7Q9beD/
FZzdcoF8ugvi5Jt6ABzSDS8jQPS4Zxlf+iMnoULXMDQDaXmwUWDLKwE+MHqZh0pF
xVUZcMaRPQyk5LBvl19+8VpIKzhXHS1K5gnmM7gBXQDrGXXKCUy00WNL0g6pZAbt
LDn8OD2RlPVxR8OFxJZuciQVg7tKUPeZz+dbIFUhG3xmnLFlczyigsKY0GxB7xUF
UFB7HOpsWV121PDhFdKWQI1w7PwjPqnP8JalSmfGRxaE4LvwcuHdNthdxzbTvWJM
SMzFiQEFahOMf5dbR95rQsgvEl0HR1n5JEbrRHMiptTfJMU3mUMiGFOSgtxnkF3Q
/9RPIfA/LGsOwxpbW7b653eTzvKAHz8loS/eDSxLZpMPoaBcQ4oBDWOKjr5Da7bw
wqrUUy9fonXMO1DcVTIafPfA+0Ixe3S4pXCk210mAgTDgpvmBq+mJxU1y4H4s8IH
gNxW+hegAuA37FRmcYdXHIcAfD+9Kx8UQz65gYD1T52Ffz52Neg9SAu+DBr06Q2c
T+5ODaZ7eLRiBwsKK+n3ks24wz223v32y7x0u+4vlKnY6dv1wq4k3/n1Bc/jKGd1
q0Xv12IxB6mnNZBqTrOBkJse/V1eloq7IgKS8aKYW5mJZLw3u7Sg63DS5BqPYx4H
pH5ZE1GqdNzeVy1BGSvy/ANa8t/oH6fMquf6ZHwz+9djK3Bjcx+lb2VxeSDzuJ5j
PQf2rMI6qCN3zW0R80EdFqQQlav1XJ9jGJF3jt/ka8KC/GIgqtiaG35JrsGsZpp5
GFNZ19gIjJz3xWIwG2tY4QZRXgSsYCbJM5II+nN4XRNiLLofle8ywEUeEEUzGZho
UYThz733i7b8b3lGuSKRHMH9mM/CI0gkcpX4mc8I4DOvGFGP4k/cMipq7wo2Gsw5
JtVgkJOinqClbX4LUi/TdER7wZFCYUk++dpjvSLU9AKUEJ7n5lbBezsb9p51qFfS
Ddxfrz5aesWZrmu+eCKCplKmqdh8yFQYH8N7L4rioVfKzjCZyrNa+w6N5O1CENK8
k+hsJTBdgB0ZUcQWlUihcTYs49zaxc54P6FcysavbcUGSWndIU4f2wlJ+xQVmq3f
WF288KvJ+vJaSdwfUXGBtrpWgodYcmHtisgzFt6JWqko3iGctBO7R93zkpKGdLJL
LAHXN5NGPPxwCVT4bCZTZjf59KM7p1LHzQe2j7qN376BWmB3/uRsYn3IN0pgfhvf
OzLRERP4yOfhefyeP11Oa48ijn5v/6b6R2SGwEfe1NBqHnUf81SGmmu7n73okioG
+wmf+o6t3xEOyF2l3LP9SG98XFWU5QtdqRGNgNc0NcLI6DB7XKviZE/NvvR7goC2
JinhDIuaV7dVocN04tlB7IkpO/rzFg53ddpk3jV0YJ/IrkGsN3VfjpOg1a45ZKWl
LjxcaRz2W8h02PBFY452VcVF25BbUIuajzpTmQVC5H7n5pvCtazhNXFpUYPnhG1H
pyWvr9Ughb92ggdQRsAiimwtwPy5HM+YfQ9pr9suQloKMvPtwjzcAtGb7uLT9y4e
at8kUEz0qsAmB7/j9xtH+CuBRv+qJbdikPXJXpUEERbnIzeuTBLvYVsqhYF5cQ/Y
5DaGkdrIRZe0HvDxmRjAMjGu9zs1nfUS44yE3JxVjQlUWKSGiUsa7zBGGhRo/RQT
1rpAolNrcOgKL4AC7XvqQm3krISeE0F4ftk9n9zmJ1Pe/XowOccxm8Kq0vzAQBAr
PyzhzhKxLkTFdR2He7OdiD4vRVAHJ/2Etw2dpTtGPrR+q2QElQdyGqAcHTmx2wrK
Khg9QyOnpdTDJhDKaGVw9NL07a9T7xy2D9Z+UCeWN61v3+y3IRLkXwNuphZtzQDR
arFy3p0QZx6UB6Io0jibqCAzp5L9WKyRGqGzpzFl9X9ixoeTrM9yXFFQOOyy8Et+
CICsOg7m7n6o3bMdWNEB9lWQr12W6vmJgJ6N7yQQH+UOq577L9P/kqXNei8qTBBt
ySI/YgbGvvGggwrLSxVeyo0WwJg0H/IbGmcCenDlFX2hAQYTSruZSfe22OyscbKZ
MKbcBB7aLq9N4nqUtcfzyntPtfg697VcAXo1k80ZqgOGnsEXoW5oDv6ah8XjXkx0
0kZsS6kiwGX28fWF7Jzu6C+uCvg9q+oaYLJ/BvK04BwHFPeoXaxHYZqk3ZjXQ/ie
/0VIiWU6tngolYqld0AUb1KvEI7Fq1gxgj0xZQdOWRFxA81SkYrwIl/IYeCMgJsT
9AEgkuizYMCq/zQbBnVm2TCwWUdKX5j70cKUg/dAj55WPNIT72YHqS9LcIqITAfm
5Xb46JF8qMBoQPnzA1siNULeu4x/xJkCdqIh6DH5OkwR4SDI/IiF9GbqCeCI0moH
pc6LhdYeBYsY5G/QNnTRDcuOHt1lyYvYzHagSiKpmB6bPXlsC1w3gn+NO0cf5F0d
1qdna+yDEGNPJcmHPzyyN24fzSWy7JP5F+h81kuOSukWR1eR14wBR96Lq72vuDCt
qwPBT8Mx8o88LSg/mbffy+0VeEKabPvUNFRxI3vWsmvdrhwugSwRsVwI8JJL+l0+
V2WDtfmwhY7YERsB+vLnyQoBPOvSe1z2VIEpbH2EzLNZWDrd0nwpqA6yBm4Am/pe
UxkKf3SP/2IzrVmfp2kSEgncnMMGFSrYRvpW6O5OiBH0LpTzOwGRFFxVi6K2LWb7
+KsKBrGUQ6u6Q28aKS1g49wb8molbfjZebeL7CFNd7aX7gYwyNHULWGPaykZlzaW
bZYL4wC3fdC+9QWxCcRXeVB1B0ZVR7ADQdTniuQaKCKKG93E41Almkf9n9FhnVOo
10T9vxOtI2jWeZ8WAXro8Oedzol2a7WX4wKlAYB5Vdo6NVdU3btbY7P6geu+QhGb
IO2L7Ie578yjETxl2Cf54qg/eDXaMzOAbkNLzHQ0g6tmqpxmLCNqHqFha+SRCHyJ
W43WwcbXeGFtcZkRpsprI7dted4IZbKF0dYt5BnJw5sH7abAxKY6t5LQFj6jlOnn
c2e4bLXzBT/IorBSxqWDVnwf765UWMQoPb+npe3tdmHe7fBad2EsTYXrOpbjOY8R
08uHQdOjosvxC3/ugdF9AUVwa7nyy4bzFvd4f8ZAGECXWjEGlljI/LH7lfhwH+Ry
UzG18UBI5JB0kiGjdgJvWgh6xtgeNAn311O8e3C/HNTvyuD1ksogTD4A5sMPAXaY
p34soHr1NxKL7qKNrvhNLk5J2ni90H28LtyTKOnnX95xN8Rdrep1CHczDP4tbsjG
xp9m4Lbmelt1DlUyUhb3vTi4m/ihDC0kLZtzuIFq69v27Ho+VDvkX0Wd1m5kBv35
gUqT7xrQaz/2+OEqzngy//oVfTQrxjdljvMX0rV7R2O03T9oC/5bF+2bzka9Im+c
nnRWPfJFT6yC0WUZAJTI8/1hkZ2hXGaJP68j7o+yYdgtqWsRLQMRDt23u62r6YMj
TdYL/BoqlucC45o4AUI3Thmm+1H/l2hpzoYQSIt8g3QckuhE+IQbkXF9tT7bVG7l
21x6spQ9amlgFeKVHUCQZ+Lnpbx5A6cNd9jUj+ZDqG2pZ8oTTF0Z5EruOD9nZ+ms
KkVPWD/1mECb4lZcNsEltRAA41lbLUj+Ue2miiXEj0EGhsyxCeIfG6f47diGO8Ee
DCq88+uL9yq//gOOflLSqt/3uyOlPgj3AmjKlvunxzBthHFsColRW0+HuLT+/JTY
yNzAIW3+4IoRFy+DERVm0vyDCk7BmAHEBVwQ8ZfLBQxXbh6kxpF8nMuHUbJ/Kbo2
wmxrGF7W4ZjAsZKuNd1Et2U+q7yVMzUlo/e5hUuiXdxjNR2hySLvmnfADYpdWlJy
KD3I5KAVuoR8ba12zsCZyxb6dcONq5yEmUT2Nh34Llgs1ZhCfm34xGc0xnIJYQY3
ZEPFM5jiYNmkAp/BFWVES4vuB1TMbvfis8ypuOJp+J+mvepkMw9aUucHs0Z+0VU4
9iO/I1OKxMEcLrMEmCCmXwumXCRJfas/asGGCvd37Q1oNGtZGjqVV2UgQHYpmUvV
nHvMECVVkR82QqG3efEprYX9Tp0BUoojjLAWu+8CEMfylDdhqIS6tGhjxSPenf53
omWu10gi/1qZOuwRPG49kPL4EHWw3QYV5hwYMFfyFRn9poRiA/6KITZ0URXCxK2n
zoRZ782KPaVhYYbgmpeFVllNtXkdD5B7IwO7Rt+KCE2rI7hjpbSZd1qG7fZC00GK
xh7knmsTZUlb+XvkzfaMlUVyhoGblikis/5sO/2KYYglQq/TdFnY8wdQl6EQA4Ea
VPMZbV5L6y/Bxks1+AeWcV4hsUZPVgquyHP221r7dJLpXUDe48voYCgu2/tjmOWb
mPxoWdIMgHWw5gv8rOIYmsTY5ttFYvWaxhSGXwO83aG87io1iaxkEl4bNtluo3Zp
xym7QXW6QLGtOh0Iu/936PgeB7v3/scovj8PJ1ex/YjHDC4Zb4EOJkfzgF1/NVNY
T5rpG31cRa+lRwm+FrhrqowKhlK3BhZI9ZkSvh8FE0iSnNYSifFNhdEZKfASWQaI
XBKOowYf9+Hb5tk1E0JVmRcbq8rcFgBFZbFQIgu1Sje7QuZsJMqpbbH2Z+8oSdGt
Vq0LqqfSmVoPv0snl03Wo/XOILNZPYpZQlL249gMnsliyHkXo2QmeB5Me7H0FkN3
kEMgt4uPXyXbzBtOMgjiLsCB5weRM+iMBJbAU2VJ9SW9uU0PvuyWy6WZA0H/jW5P
FIswiyOP3okneca6h5WsbHZ3dDFXZBKJlZcSJDTIEwhmt8rb4WujQEZP75i6EZzD
ia6aVu3wh3x6oWBCyoHZzGljkRlQVWVsv+fv7nYCCIrY/h8YtCGBU7XdzElxSh1n
SzAnAbvCN8ap7mdEBc56Orps+BV2PXpjT/HwZrfoj9D3w2hTeaSq41YRKRrtL0sl
uVc4awE+8+BTEbB98d3bUs5aiqOh0ZMB+wyK9c9YoLaTIKVpl4aVkACidxrOCTXG
9hFsiXDTz3TF4IX8AdmAhE7Pw24c/2+mT87/WGsAmlZ6Ku6GZxnGhn8RaP7IAqju
cESDP1Emt0AyMXtDU7JQ4GDmIsG3r1iABYdRVjo++kigPxdsnGP8HvIHFIoztNvr
M6UZTy/+FZ/u5WRtLY43YjKgzsMiqW3PQg94Ex6TP3dOG1Fyf7AZ9i7J9vIr0ev+
I2YKsLChvFm77SqjS1L3f5C0kSBu/eSCrVaOrRoW5neaNZTgTpqgx6ga9Fwj0wzS
jB4LuZgNzr4vE0RLdmAcSPO90brV+qc832j5tiOU2GVfj/XNwbcYDqp+cHNzl8xI
0+XG0/9Po2+9gCCroUTXJCOBxhMCI6IbuDokSA++0dICHSLBhe7lWFSNYFJpvkuB
sGzFCe2s2AzEhUxFFga0btz7usi3WvYLa5FWzbxIdDxs+kyyQc4InEjiPH9pE1qN
Zj/mm7+C26cbCJFodB9bLkFnWJ9l2AEgtzPQCUqtA1ZC7LIuDEWb1XYefQgaQo/Z
LvOTatnQGBUu/1T9yTLLN6q0Xv7qm0qZo3mCok8Q+DWxtg6ZRN/Sx7euMULJ/KK0
OMuHr6vSnPDY+aTM/ivX4s9cv/KKL0KQyDYZ04wJQKQwz/CWRZ8KLSQf+D9dHDn0
qN9rOeMf9CbSnpXD4RmcyC/Z68KAQPHTqEv/3EHgECsHRR+hK3Wjdnk4k73hKiNG
8PQgVdDdrb+YdHWupxn0l1jmAUGhqT3lf7AZsjQCeA8Wg1Os8KsaJijgztxf1WTE
6GkHiMlKfvPBUCY81FeklCRuKSsWd82HBKyW+N+r80w2vdp141M9SoQ6JC2V37nu
ldiodsbLIICzyclB31ZldQq3mjCn3obDMQ5lf7aOvIFhr1HNUSrPm+yAOY7Gaqnc
va9MNKCxMQALDl9D3dNAJHtBWjbLSRGK7wMUu8cW1V5lW6JezlrwRcLLXf2gII3M
C/gm8s7ajv2Jvpw43lEQEnHUG89Ve7n9Yea+3mqfHh6lr4Q5VtKJpHRIXBvPLnLr
lBvMQ3QQrFxXxsQ/j540o3tRTJ9kB26HQ41IZBXbwsNS4CUImVYkAlRBV6EaZMJG
w8ycqwD3tdnijvNCkSSn6PT20+YPt+1RiQg/NHUiVBI63XJqKcxx8OZBJb2U4Kx9
tpQeYolNTNdn2h0EqA5tJCHJELUUIHWm/DeRevTxNS/CFGrSVZ0Y2yeaYJnCXZSN
5Pndb/T68PlaF5vRIshftkw6g5qpWMGqeB4VgLXji6r5aD6fPzk/glsqbNAQLysl
0KevIo5MbZHi6z/R6WMzTp2iQjBqQSIGfhPhnBwRIreGgnByn6G+6JfgNvPP+zkC
MF5m5tR/bwuVu5TI6UQHex8t4QTdqgOeTxWDkV9AoE86xKJ9JUiVrnu2G+F/4JA8
pHrx0hRjuGrG9HqOF93zGnRSshjvgLJWqr+iQc2N9vEFtNz0AASgxjRHu/VBdmWN
sIg92IzZ6cDQjloB8HmTblFoM7Z9rRycfu0XmNY7ZX3JF+9rEi+YqqZ8AjR5jyFB
x94jstRraWBrrRzOyU58qtuEsm8LgCTp+FLBK7lrwszsa/oXrrpnctutoBKual1P
7z7LQUw70p9PZ0R4snx7QIs/43otP6gKR0hoS9OOOf+/k124w6Hia+CoG9UIFJHo
aMuHG2MTd9MvZ9pHWQYEbIadG0XH72viySC6uO9tI4IaAtGSbgkqwgK/EuaS/VPE
9E5/IkYC9y4TbpW1T13y8n/C4B+W9m14EBIIfGB0uNrckV8FZBHlOheCipHUZ5nZ
066TgWSc0pYrVe1ys/qK7D1Yz+kLZymb7vAsJYWU8d5jbIvzC+PUTo6cd46dMLJQ
H8gjpBIFKtE0uLLOqpI/IPRh9vPwDa1lPm43oBXkyQIo/8LyCVSUsDHhHF942Jl6
EOodJXWQI3oBTdQPSGMJb2L/a/wKbVf/WINg3HYSOk4kGmW5RLu8bzyXBMZ8YB56
7JTUhE0VU0aXvxC9LXTVveLoV3YugACHxdtBggjpKZ+3bfnaFjB4Jzw+pkhCWscp
pkXb3OTyvjEjJGnf1yVwC6wGMwYrYLF+EBLmNijKshFFyzdN/rThbWuTQTdMUhld
gC0b/RYEG+AXnZcCbTRIzoqouTeq0FB5mMt1JkkOTS6UUIk8XwBJt2bKnLxn4mD0
CeoxIDL4IsOQDauQYsrILBCjND/1YvaSA63HERQyYzvDm8mKgkNrpazzqh3/ru4f
NUueu/YAE1LIpHCAem6KDFFHju/N5SVyx2EreHQP5d28o/GHd7cvDerqKObsZ3pK
TgUgosV+EX+wtjun4gX54Ajb5NKvnNaU+L5et1UZX7jV6aJC4O64dnX+7LqYZ6jB
/eXDMoOMe4RgCJ6vkz5gBrjs4wf9CEsJXR1OKNmGCfIlYv7BzumuYDK8CLC3EEXP
wHTQvqeNh/3CEjMLCODdqHdsilrvWuzY6N9M7xgo6CR6I/9d+IhQiy2LGWrh1OAJ
5jM139/oatF5GB4fHmFEdAcoSbUXQJ5MDoqiZQ25AeS2Fg9ApQn8La7l0aT15aDr
Tmdv8rlLO7LN9DiQSztoBb1/RSm2YYPQnRLNZjyUeUj+OeekPJnPklya5Lefqaj+
+uF8SJ3shYIp0BPCg52f7evEcMUXEznBQSY8hmhkX9oG78RlgF1t7T/tx4Y+jTfT
8k7keXwDfd8n2K/oTBhUhRRkGaGvv9Ewwo/ve4Z46yCYskSKn9cO64LCBkksbYW4
CT3fdFy3lSi0Hev4B4Fvzg7/81AW+MltMjVptpFFfMw13lRx5rfqM+0wd/nfeZC6
p3bVLgjRhsHlzLZ3B+lZFTLN1VmTzJd6qlOd3fsIxK76COMFdznZflYSHVUpmOgO
fcUJBaoHiBPASj12zI0WBucc4hMXHfoEmX7qxhRvhfxP2EqHtyDuSW9Xpr3qW4cf
RJoRtQJ79mwBsa28tFUh1VOTmhvMk78IbTej4CG2hnzifqTYVsCSSlnLFcjYU8Sx
ANZ5fLup+4fCuo7B27d+dqIbekLYKzv2kwvh/tirk72imJJkK4Q4tcELoa+Rfr1z
FdKXRWgjAZJuOtv/IrEmHTX7Xr0srfEViHL7DgN2193bqEeufVmtYzF2kur5BerC
+T1nDd4pGkLuiWbFTqijnJRewyBmQxXZh5d6d750HSEZkCt4MlLBVI9mng6x7mk8
fhWokMoqcE72eXVZtcguinXatsGqvupRz3OYVg9PnYi6eMv7M4ebq/xCx89sxLON
Mkw3s744zV+6oq9nG+O74Pyf5ekUWXgkoP4U9WJni1oo5OORqUCMZi9CSoCrmOa1
i6yCcCyA2eIOhu7tU8mK+oCSKNJ28m+o1jxVjxvhYPvBAt9Mbw8m5ByZEI9Xr9H8
RUzHGxOyisJ3fsn1QOm/k22hXchZUBV4NGCnCwRjRiNvzuX9gBLX8tu1KXfpgJZy
bwspSVDj1EE4BpNo7a4Rb5G1HtuLfdsR9ayA9pVwzTrwGYjgzcagZ651VtDrk7wF
QaxKzR4VAmmA0AOoCPzWKbQnmweWEK7HJGoNnI7zuDEIerS+j5zV6pxQmTu7XsvH
onFn0/ODLL7gDIPjvnxOkMX8ZIH4UU3blqo3N8jGgNdZhOzxRQE+UYGx1MCWtAkS
HSJBhdDzpHQafmjSLcFCsvgP819Vqi9JeoyxfAoqclU0ueNaxUw00NGZYYx81UTS
T04Nae3DtOxWbT9zcpYxauY2UCPX2kNIvC1/lVjxnYE3rNjA8j9TaW00aXqW0aDl
1LOscsIKVgafTpdPNO+J36Dxm1u5yYHg58DY5ZShmXh8OV3/Ws8NklMzDDYtjgwo
dkUiUaeSllnudJQVTTTbHjaRbjHEg0vJm3Agpw+Isdr1k8mG3mNZGpKqxPRH3onN
SlCNCHkw8B65A13d/lfxJ/K+4KuzlgkzT4/iSvc7x9biQV2lokXCkqoWTEhJ7UbU
njETJah2cCBfpM8S50Ba/ha9+taizhhsrGjWXBg/LESPwTuxr29IMAUE5C01df1J
MoKZs2VIcvrH9mZe8ZwhjepHrFAXNNU40tib1dob4u1pKKLUcGLqnvQaSAgooURH
YEfRIK9gAz4kEYKk6Ok/5qiSAEPOUYrQ7aQhLqskd1L+priYLhb2xxedGjQIWUt1
4bb4d2njDdJYgJZQonVgXSkr5p/Iumo186QWNPIbeR6xZL593U1c4x1SnGKdhnDg
EMnloeLuaTNk1aJGqV/jbhmzz84w/nNkWbFjwD9q8aT+sowWCwRpc9n3bcsFGDMD
rWfq5duvt+pyVEN04fqTXp/TvvQ/yBoN9cMRrlUZyaMa1wkoxzKKqTAwJbMiegrz
gunXNuAbBzPSScDdd/hNq2XvMzStd7IDC8FTgjVEF2ZTL5Vf8IrcvEyJ+A9m4tpZ
oEPIj5i6qQB9BK28xGR2/u8YX8LMHCdpi87TfU1GfienJ5GcscH78kljT7MePH/R
wsa1wu3Vxv1aC3omm5di8fIy401ISPueM3EoCNqJe9nB1eu5XT+NOhB/47Q4jHhA
zCR9qq/rCYHKpjWacHQPm5gAt5E12ZOJLePKyNYpwcZL5yJ2aKuIH3yBqd/3K+Ca
xIG0osN/va80KxSlwuQToeMFqF5EbS4tullgjFnhsX7xqDioS9naO+VOavesHXxj
o0seA1lTZ4AnzHDHxOC5HtnyDe/Uf/QSud/9gTR3luzsyysdi15dvrjoHgBU1uoM
SjjxbtQ7PEyPw9uRSI2eFiA22lh6XYvsL66A9Nf8k2YLcu6mbSCA6Cfw7wesYFrW
4s+GaEZUYzCOMrXZBi5zP0hNlurerkJZrx8HkgT2XKm5Q6QyXupN9KraDOx/CQNy
p8LSlMCtQ+q/EIAZqR1m3NvFy/LhHjBDXW8r4LcgyVaws2rbS7iEJ016KODX4y8i
+0zz7m3aE9WpFEAlEEEt0z1ZGUDG6V/RVdc2pBT+HoHemXBJACefwnFf7x57tyOq
xmZxGHO9zDu6nHuPBAO9qbTpgC9PsggDYzpYz4b+Xa8j9AcFDEphCo0xHpdC1ZA+
oMfXNLY5iIe77TsUln79VXMHV1bWegZMvrb62FjeT75Aa0rqPORlMw/9H0iTJ/yu
/f2frTdSuJFrh4ndFWb/v7/FeDNs3sfOk28oCWCQR657bLjK3Y99nw2tUmUM/VLl
IYjHJr3DM0wduyrUrlb0daQy/lMBMELNUDtEECmNH8ekzSDNR/20oxtoKK2bHIk3
3cR4EeWcmwonPcWf7RKypll6ctK3+r0iEsKPFXeEw9kTxLVTIdIGNupvtJsHdjj2
GJpD/AbCUxpf1MMdfWbGD6jW/4b2foiCTgj5PaERyKI7wQZMzjqJeTxTKq54KVpj
N3VjW8B8NxJMi8b6KkMnIG85/xrsIf2mesBvV09L+yD0JdCYpfl6MQxWzIcwfQtg
sNfQ/nVj786VaCCN862ZhDM3X9Qr6vse8NAvK1GVjQSt8QawkS0x4O+y5UEY3+Rw
09enJjSLYZYF4/CQwcKBuYvruCSB25bzYKBAMo+134iACdW9H6IKcymNV6AkCaoK
CNwg4E17N2YQME9x3JLqZgkwKdyeOKlvY/SN4KDXY07KQVwSjGQO1A/8+72PVD/s
gxmWr54EOZ1HZ8xKhFcRLk1kQ1rc2LXiuvVbyasvuNAS0HtTKMROqZ3zrE3S30SH
zpRjqTmS7TRbgWbvojGhGQaAFVkWZ/0DpKGvEM7kaqEw2uEAlQ6a8oa9vJNY8pYR
76UoWipidXKggbKoM+ok0tma/7nXVDcQEm6Wto2qaDKgBMoMOmG4sgXbXhMQd5s8
ZW7t2z5w7VGC4CYqmsXUHtSy5DgyQ7z7iNSyTlm4CB7t021n+REYs7PV35XefmDb
lNO9//cFKP4J2F2nJpbeGuLx0Jo1mj7UxomtiafjQl6AS2rf1PqNLMHfYqAS/4Ip
5SrkihdDhQcx2W6mNjng3G5HoDYQ9LeCJU2+K7/xxzuZiigNO6cOfxOO2gNRE/SO
FKl1PRamBQRXzBUbSikQB6BqT1K6KKN0PsvmjYt9VOHMM/Cbp/JgfUTM/e0FTj4M
v6wh/J67CuIVn1ECF59wMX1YRu9DXEkYdJzuqo7vxh9QOzS37SwsOr38v0vZpyVB
F0eZiZtiaZlGrei9Jf+DeOE4bM9je07dZdh3pP0Y3kiE8vfperUda/K2PD+QHyDk
lq8KJqB97JmmXiCmKNTQNVafdlbk0f/Q2bn8o8I1r+Xbi9KK7yJr6ItL6hL9Q9+R
hOHAZRMqevaeAPm7TDwEVzBUUhPR6cYKbO8lNIP21+NloE36CvJ5Y31Xysqv81ii
i7T70v8+dqXJfv+nHTryzvgUiWi3k2HxMG535yruE5YrjsFJl6hrFjbr+ueAHvGp
zmhFeaNUwUqvZJJeDMZzQjoR0WhWkn1pJfmWpEXo2YpWob5w5y4Iie8WIFQSkP6J
WYGQh4Zp7kx6/5nTZ4bCteHaB93yLTIu2i2PqNq+OfxGB+dR6PaIJwx+fyedwqAc
NMRhLiIeXtMDIuBHwJoewewgBUhedLbMy//tF6gHEXP2tkgLRrntwsptFxAGGXqC
kYxHlBzDaxOcpgjT0iUuRmbZfd6AE4K1CRr0T1dFwxW0Wf08KY4k6ACdqellpxUQ
XIWnqe5TJr7QDDXyRvGNEQS4uOIwAkhhnb6ePWyNI/RorZ1fkh/BKmnwugNide+/
I66WzrKx2grU36FnNnWlGfuEmXXCpj7t+vGhoI5VebaD1ipsxJY3PaxkYHLxuZwC
uUPgIbw851AAYpe4N8tnXVz0wIcSATsfRzw2+4XLTsuRuLQtaR0TWbTuOIEDSMUF
CuyxMTj9Sn0H6g87LfcOawo6ff3JdUAkRWQPBCRrNAQ+IJcWnMVrp2FaI+w20wnx
brTiqgUkLtuMIFONuVZj/Kec8UjfIcAX5bxQ5z8Jq9jUTJzm0Bzae+8lxRlsrvYM
Ekpi3J+LlUOezecnWcgN1LJhYnoomd2xZa6Rgyea4EoyAV+ibYjAv69Kued5rfDo
BgrB2kmSI0GqrQsSc+jG4Ca1xmgZawG04e/OYbtsPn31hYYKLlqEXwBIw/4xgQCj
8KrHgHFtuy3Yh9vnolEPwyrUej2vFizpe8eQUNYmZaqqNdi17d3/mOWXs3CwT3Us
uClsx2bSyLTYNBVng57OAfJb1fnRg33xDdM0LJsHOIQeGmgN9hdVa919swI19v/y
eP0uwh89Y5prsHNoeZwcKpuSJIRQM1XKoE5fE92z3YFd6wVwkRk/B69zWnv4nT+J
o/obLeuz3JiRaPQUkVC8D9/r64WAp41uZC0QhhoovMZOQ+kWyfAd57MUtOQ6lSCT
G8ZSgCiDk6+tVLxZNMbZ04zn38E57xxsGOHo8t2k/cZ5yTSw7HH2xGef48jpRO1B
uodlgMOpop2NjqqZcpEJMsdtHqKnhXH6ynibWJJ4YmKLrqW+qVtjyF/0n8LcQB8r
jS22Do6ax5jcDYAabmKcHWjVx+O/unGJIaguXD5F+FHfFCQC7GhoECOjVD31r9qX
1DcsuZHWb1W0fJsZxpbCdVKW8RwD+OuJqnYH9ab+XDPagC1k6NEY9BiVJKX4juxW
jPO7WH8OKTtjPwJv9e/hX/11Gv+JfuU5NNy5YQBkjCioQpitSl4WaNJgZM1yr7sK
pcQSeoR4DX6Ylu+hV2bP08lvrJpymQp2julun5OzC32ln/wlgKjcfnqXRMyF6Tux
wOVAAZrf9lShDDQouIJydkjBgK9csKm8R2OSBtcnTq4xKWhTDvOEF+GGj96iURm8
tfWV38h3B1FAa94+qUH4Ouu741/DobtvyQt0zvQXdhfM6maO6STKNrx+AV361Q1D
Wrvw6cEGX+1+TCnjLGhUmyk9aCX3rn2eEKfqe0o7KO98jZPsnd5HA7FuJwMz6jXn
CAt4KciKNwwTtKsZc6DL6vmRf4QwAhYLsE2EGerSZdJkPkLo4edus+Yg5YjpzXja
gljWwwlJIRUFOYXrTcYGFuOftPOA/t5t2iA0z7gKGZutBarGvOiQfk59BtWrwXHJ
krnmHprUOx+InPrb9PjW3Cxqfi58BJGGxUBpPGOVplmjaQavp0VHi5V1AIZp+zSM
OxhQ2xQ5Cd6TsJRNF6CRtp65k6yIVqC4CIDvCmKFTBJAYxm++ixQHUxKTzmks7iv
W/bwYtcL6IY4fOkM+ZnUWfbAI6d7nGnATrt81CvsaQy/+Jm+D9fZFpKDl09Gp574
5q3IHN7wz47twN9hzcypDQYhvoPaZJZhbo5+m0JdoAgGGmTYYo5+3VK9SzetUZZX
tmz+LboEEDa4lHFwTlIAL2qSpTpknby+pPRpL2ySNaI2aA/u6BLozaaiFZAamIyO
KLU+a0ySRizlUKjZ7liaCRvihOIznGD3zg2Fq+s+GbZ4j2AiNR9WDuJZocY5RAZO
eoNGZozRajjwsDMYgMUpgp2UvtxjH/p9kQ+8K49zsssAUvUJKaXl8EGqJ3hXEyku
BrSibSCzFS3/QXPqlgM4BNfBLaxI4WY6rMnCOsY5NgvKjVNIfab8eEo+CVLVNxUO
ZCA/QpMGnJ2ieQ6NS3yPffmYtLraxst36+PBEFKDqQ2HQa5QTaIiK1wYLj5MKw1S
ixNR42gB84L4NfuLG9VIRnl1ZNSD6oQn67sj6dqR/RBszfTlk2/tgax13PsQAyDq
Gkvf+GFgEBZDZm20Kq4lDAQgXD+2INUJRTk+LJ8HZNoB8tanEE4QzibbUqV1fV+l
OSHics0NP1bSb9VjOvY6Xqo3EMKqjRK6s3N+plZsy8QejfcSiIDhr5uDDUWriDgi
upjBBoaUdqnRGOPKac0u7C9x3vFMYVxddzleU34px6RXyxAkLoJd84lB4lepLXHj
9lkggIuS4Z2PTPxlVy1USDO1N0gNC34QyN9N8iCZ6FaBmjOErVGc+9W6nHPrQC/b
Aqn1O8dnsZkgFuc77ZYwF1ENvAw/kwzQQ/WqAeqFySvP9mzXyov0Cy2/gPR1A2pd
ijpvoMGpShcupVH4HOmOUVnfKdgmticC/D0tZkQh3i9bHMnriU9Uftp9gWJAqOFk
djP08V4/P+l+OtI55VHUq7ake5QQUNfHEuBquz4qhpF/j5ieGbdi5PbVOxi3XtNw
1v3EDG91P3dJqxJYaUGcV277ZL6YKrXJNNGidLCIHyuk8p3wlHBBbIxkpnAJH7H7
m4KmeGikDHRAofgE2tiwvLYUOE/3pwpxd8rdhwD2M0A0OYNpi0bOHFXLNZXScIWM
cgOhyH9rrPoFAOhjJBYhFcW5kxrGQVQlqdBmMytnjjNsf69qgn8v7yRQteLVTVi9
YFfVBZJMeJApL5boV52999jmUzDmFkP86n3DPuNRm3smCNqn14UupCZbcSSqPu9P
UZsGlyhKR500fkMfu9PI/vCREZzV86Ot6Onco1JTBX4+EWwiFKCfVHt+dCz3D3P+
2B3oHKpaZK72c00OokLxP2BMvO6HvndnXNroSq/hfpTD+MJvBUtxvvcDvoA5id/i
N3WWHfFOKqXueo5WKKsJ/Yf+81MYsQYIAuLzgixXipCwE0sAZ8wwcwdJPP0uQ3/m
Uw4cYS0kRCnyYLrx04u7alBQVd20i1ulT0d6EKWM8gi3pqIJRtB/+DBSFATQrwnZ
Fe9Q77+wjuGx3HZ0L/1Emqc/y8Y4CrOiuCI9nVzk7JxFs0vChwStn0LMK0hsWJa2
rRj4Ft6NHlBZS/NQg7QhjElToc4r02QuM7FkW1tsiukMcKXX59fsO9Kp3lPYFZC4
Rn3LKuf8+qLqWr6fBhtRbjYfkVcF0OHI2yy1EEtIAklebjV8Pp+oYPZHHclNU+bC
E6DASzwjAsXUpemn5bLya2PkfDlX+81Q+iIvZG8Wx6v/MKRImJBs80GHbMfy2Aua
sRVB4SWpdcvxK+ETZfjVcUHeGReO+98eD9aAzs00DufLroB7zl9YNXi+CT1/dIem
gGOBVh5tI+Ki2wvI8tRfDpmcr5LM+I8ycvkLeBDbDJYc5xQZpyEKJl4CY4tRCrah
JqDYxBDzezfMVewCpEtOtuglJIzOsYF/Jbe4MzxNtpb5153AmKcTn+esFAVWEspt
bt4st23fuAwQ/CT+SA9J6GHpHSE1UdX9B1lBVrgR1GgJQlc7foTX1L0xYRhNzRp8
YAkCjORmGO6GM12cyqHCdPGK64lY8zyYkxRPnCcmqzbyw636To4GCHdOa9JZl8CE
QHlwC04cbja633XdZjX6pl4Yx+vB4bOsazVrKFVeKucf1op4SafOm8pm8VsNGC33
AmcYXMnaCt963jWCaufpv+PSNwB5JIauUcCEeIkKvnVt17vtD04Mkgx7TRGBFLUF
Hrvam8q+jEGmf4zh8QBrbpZsBl/BPDG7b3wfkTd/oB8Nmk448gOMnsnWc90U5pkO
qXy+SN6SFMulyARUw9PGVLxrgHSe1V/6TrYlKct4kno6YO6iWA0DNBzNZ7iP8YCa
bohcsbyFcFABqeQSN4oucr0k2CgY+8k3uIFua/EPsoTGiQpKejyeo95yiazw9mUc
C5X7jsmWvgU9NgxbPzvnMjgSyyBBEswSj2CGggzmikjC5LLplJTPk7VNvchFoAN5
O/Wh7TdfIYd660cQ8irBLn9bLeuB8jBbakzWd2fg9qNKs/uZun2WPyV/bm0zRDgE
unso9HQA83H9XJsTZkXwQVDPttNZGdbq2Ht1/ROYjRRUBJ+7Meu908F12285sb8z
2WGUFilAQwB/RAcPOloEzvXYHsV+5ssANl/3O4RMgC0G/Q2/l0A1p03zE+Wa1mn8
Pro1vne8sOjMGTm3KXxSHR+qofyNpLnrBqmh3eg8+jS8xLNwd096a6my2r0mb7jV
qk+HtvrjjRTHJ8vcgxgCfxGCJ3KqpPmCG9ZdXSsoWF+JzoKLbt9QKzm5Frqg3TFk
N6zKbNm4BqoV0ZrtNxYnTesVkpE5+3gtyRit8sdLn1Wmic7vE++Yygcbvxvk3r7d
sG0egSYme75gYqnELTs7Di4LsH1tN7XJRV2km+F/e0a8/5LHFw0ElVVaFzYPfPc6
8O/wDRMxbTacCcsjf1DNc3STG3JwRr4Sh+L+JWBW+iEMOfBi6ps1Uo0ELtLj58Tm
ZvfUkOw+/IAPDIH5l9cqozAznvf1PdV73+Wbveund1eBmxIT/49KeTVo5WzyLB7w
44wbVO1NfZ88e94HhXndIKi6TrZB2nsG6d9EX9LlaWFTp8ymY38nEHm7ACG43IcP
9TWoa8Cm0Ad9GhtmcyqLjmZeVWddQFlU59H4VaJwCzx/bUMS3w6jdUsxDMyAoM74
rY8CtGScb7NnFBbm6s4yYjZ+KNRE+tsZ4MEZycag99XKXnRluOIPYa4jwQi1WJTy
meyk40hGIAXt+6AbE7mD7dPAv/bTmYNOj4CmyfBzGdH3s9QkWaMeURceUt52iLGw
ZjUvdGcQJh+DeOywxgU6K3CCsohrrw9r0QE/lUPNIyxnvteDDVIbLszPr3emh2/5
jIVTLovM1ZTX4p2NxO3EbIHVf/BU/VVfZEAcZa+V38L9sYLMSYYLinYbsKZCDewd
RYTAwGWKlgLbQ/kI3M/mseRPN7ZI/3TsizrywF3ZPkRIwLOCKrh3fT5CthHHgKMm
K/wzztHcbeI1WuCnRccTNX0AkA5rKbjPRneoBMrhI7ZgQLirDx6JMDgcWpQbZ0sR
hVGui18ByWxhlLAMgpG0Kxj+uXBcvz92LUs+8f3taAzUQiMf2v9LXJuZEAbqCyF3
Pz9iEjI27nmNlXlYPKnwepfcH9qsqWXgxorsZ9zwlCrVngbhmC6TpuURZYS3HsiS
EHNnZH6qgCVjhlZWq8nI4j8pFpdhsH0BYPl1uF6ZOBR1NkJbCAz4y9gnfh5q15W6
d8zOgTHXvTZ5Mkej/aqXkFrpTIFkqnCKB2So5p2Rz2/3awNCDLapWfc87TaoT5lb
hXeBcxaYEFX5+g1iLpDEByAicoDEWiJ/RcgipZ7z6d1hNXouX3HIoWRh/91EgWLf
UBI7S9ngEOHjpbBbUHnEd5brU+QtH/kBhhpAXvW0uF1qDP+Tu2QIUmw1ImUR/qDj
uLUlnJkui/P2YyO3NyCGdsac7UPInMPC6kuGMga4T9qqeno/IcxuMxx4T7ZLeIAx
yXdfur0oYLDaIrMrJdj1C7gZw2OtJxDz8wItTGxpDxYwo99Gja2mAoFVqQuIV996
IwgzPJWx0TwnorI/PFOA2St7LGCix0X2hn9YCsF3a531v2z7uAVhBA4iRXzXGgHl
RsGAo7LbueOoxNzGVdkswiEcAWT8bsAUEzGXy3AkgzU7IjBXpwM31IkaGRS8g0uu
NabWlQ+E5s1niC19+zAm6w9hwFF4hqCvg7Bvrs+iz5TDL/u23QaY3EDVlgSac7m5
/BIWZZEgjUFqRnPac3ELXpjIouYqyKBpymgZFYdiIn1mYUfXV1UydWMESj5kyR+x
chYkS7ryGrtpHwXPmQ7YqGC0phHSLy3tiXHXKwzaO4gE6tkCafdJfEPVKOh5p6f6
KNenKq49Bs0mC7dfd5GjYYmMknQuoJ+4QLdDPnhoBWMSFIe5o3EWKtAM0k2cgiKz
//3hkynn6hIq2vf6OwmnFFSNwIit/HLL1SLCskqvXUs91QH8D7ELY5QaMwE7X4GN
LgQ790PfKoEElVjHasqc1whol923l0812agPxDluiOwyjNr+A8TYZ/SaHfIlE03k
+nMLPhCLh4PZAW8paEe/BEnDXv1WpPfC5bWWv/iWzrmxdsiNuLm0f42FoSGGpjkl
W3kIGHDyVOHtInXFdrQ0OWjuWHLylftzatzfq8uBJKF3Xm5autgwex87iOol0IAO
6CoC6LXkaFH3/tU/LNYMRA4MSTJS93nM28eOaWtCRxDQz0Af/eXHbaaX+kdxJg3n
hFC8LHfuaSoyHPhkx8yyauxG044v1+pjse6je0G8dHHj0QO3QFynHjs9sPZWlYAw
pN/zWs8snx0pH2lYOWY9MfFRtE6iuluKYcIz04zUVaPhBlLReTB85MtAgCrZB85q
GPxx32hlY3whG2m/owDOudaQvTgFXqDdeMinTICmzuwTlpdFZoXjhfoDGlSC2apw
SFUKgET+YQW/FBHvvaBneAbHQ6WVvT/3YybHWUDc5M8h8pc+rIVp+RsPfLzO/mGQ
TBAdzdXoX3J4B+Ccm7S9dJpZy7Qb3JhZ2zbVXu+kMdIQltkBYf+eYt0TH2AsQF3I
EbY8b8FxJ+PWu4x8QVI+LtNibdmwVEUbbkOPf8GCkreb5dRZPjK3fhhwKw/Za9uO
ExtBIuhRHxCzW8wjoUgTOPRn7zuAI6LKJoZX0tOPjhb/BYeWjKZ+Ji6FtN5sKcan
T9QWEVveJUD3rUL/8yhMFGslOy/h9WrVYqHpu2y5TpKcitHppiy8+OIeJWoK+MCi
eSCk34LpU+9Mq3zaQmvvq1hWPj+gwoOHiPOTjDJs/313zWN27fZ+kkLGsveyG+zT
LCoii56R/uXceKzu8NSYBtcmAv/g6xdK4QW3/WWVwBuLljquCCu95DdwyuP8jZD/
+nX6UPG7M8uG6E+VWgAzBS5mecJUobpnPK5TA1it/N3PUI9w39PY5rqIiqi7N/sb
Q8dhetvroyZ5XFr/XZ5u+AP1lPCVBDMj3yt2jPVuLZ9X3JiQ+pdr6wsTIH15HvjC
Ulb2a9h8WYDOfz9zz6OVBbp7TyVa/pX9HOKG5382ZfTlyM6hWUhVHKEAygMj15OF
xmcf+24ZnuuqIdXXe3khNetb2wBqMvx7AlF2zqGx1ZJzoxm8Y/n95OyjqIICnxYQ
F+JYHIcCtPseFL0qjz5tVr/2JWePmNtnnFgD1qxyBtcwju76DW6Ta3ONhG2ZsSgG
ZoDVaTiEKxmuqn7WJD2xmpFpGrkmlZlQ48vnmEAaRHWF9q2i8gzDIBCStDty/ybk
RXhXO4kkPz1Kte29izHj1lWepGpcYPcKqzIrs09bxYod2jMjz/6+cq1pTkqPuH4b
P2BafI031OlSuzVYGae02Rb3hPfpyLp3BXnnXqQe4RT08F4hhJNZlD8UZyUsmIuc
qXVu0VHMNaFYGGX0mavw5CSphfMdvKEC6IMTXO/DEPKeP9mM6qIxmJQ09fcGFlpM
rZyoDN8QT4uDYzKfRCRktTam2eQVsI0K6s+nVN9CLTmfwFR9fohTRq3g8rPVs2ZL
K+s7ShL+SMuokTYTAB3cVXrfPBS/MT5XTv881belEJlBGZCoMDmJaeEvWXbBXPnP
CWpFLlRuUxkYkWfezJRlg8qZNAIUyT2yKXpsdYFM5MOA0WA4rwns3uLhQo2worsW
Gt7CMwmHMR6JcMVST45G223vEpYBuyW8xMLkLIVyF3ouSTlNS/O85qR7pWDU6O2X
mTlc7XxxK187DfL5HYiWPV7GiHtMqgx67WLr4QqgPUEGQpCRTtC7xSKzmowQt9NW
ONwgT5CVVwtHEuLUpC3IAIVZw+F2/eYq5Keejr01pT6ITyHrb5oFV/vhtivuVZH2
7lRTlAM7h3IHVEITR91oHOzJPdc1O2yTCxMI0PTkmZDbcyx91UD/0jI1uY+VsUKa
hlViznJAGKuM5mxFELac9w414ukSudXZRvnoSnTntmOQHblpfw/40XDCNdFD+l5R
b30bJhDJpTXUNaPv2eYU3nSBx+kA8LPzzj0CGQLHJ3aSGo4xiJE7maAlQoX8hCLf
YoOSMYXcc81DdyMpz1Z23kq0gI8/cwRuxm642YWLIe7KouTUjziedMdIFbULcycY
FOhlQldYaw4lmrUdE6msZIB9Mi1aHfqX/f+uPyh8mKQzUHr8fh9DcYVknpbeVHYa
CkkQQeW0Ea3avxBWwoGigG11FVP6ZE3bWh0+Y4ckwJbTvAGm8yUSemhA/DJ/aJo5
KCHsx84K5idNuuiRmN+lIMjYyVB3LKpQhEq59y5rOn+zP13YxbmeJLX75XMgJmVN
J8Iywobd21Et40m+f656SMKEU/6iptsfIeLkES0e02xRh3dc+3qmuCMJY1tJsXxD
WHeV4Gtt235B8LaRl/kBcEfeAwgWM7nAbfg3YrH/ENn2qmhSmiNrTyW4WDIF8hTo
y3p8tuQmhd16m+EZUBdd/hnhlkP2aQ7p4L/KvkvGMK+aAjufbqOOBHQfzKMfo8Jy
FELGPhtPwCjPw/HiW0+KIZx6JPCLNZON2Lk+PbxzywanwSZSTd2vCcCT9KQ7wSc5
xFJm3x6skMUpOOkB0uRdyRCO5uGEE80uREgch36er3XAYUrT28W/xauT6peCaW36
mN+RVxKsomlRwm/DkX7Xx2WsR/3z4oxek9L51uedhfYvWYxtjAzL+dlcVhEc+oeg
QCT2STFYfn7sabVO6h51Kc1HfDlqzSjOhHdjHFmaXFP3687AaR3hdk5VZx5XAMOg
DATufWvQb0J2bS+CKV1EbjNuH4och1PjK2e6/S1o06x7eLIsuRIOrtwyUqa7nydF
KvWbGJDed4Bpo4MB0Xgg6uqo1C1wj/T8HgStN6WfGExjH8jl8cjIvt6+pnPCLAzw
X5+TqbuI+L5BKZYmrARBVEG2cBU4Tis236T7F01Ktqbwc7LyzR+kmkcrOeI9Rpdd
l2UEkhRUKTg5Mb1OXwwSONWazcAdb0HQ2q5G/FAUSZWbYJgOexW0junQ6QMvt34p
13cMjMI9yvBh18nhuFlFoR7XO4Vk18hV7SSKwsx0p78QEqT21c+NLY2oshttncnm
l9v8LQH3xgCxC/qejcogYPl/wxUk5OGSK7/sX/UYrGUJXCtFtA2JyTHNm/qDmOp3
tMxI4b0jfrTIzyq0ZTifaSaGubKHwMOftZ2pTxcaAUvqSbZsBTBGhi4GX/tLjKPg
9IJCxb9sIZI6OK6pyjtEqBCtXplFI5We6DNrlBlsgGghD4I4UuYTlbI6RMe3lsDi
Whrx7/zPC27gFAfmkCz+bfFBNrMFBlaZawZ38Kblkgdh4vyTibw9rbFKY8MFMf7A
0Fs3O/ARYbY6AlMZVfVHFBEvrYmfUM+NYLi+KPRwdfT++U+t0oRxZ5P22WdPuyrF
dxe7/vLEU3WDf/vdLCTuSCqWWwq1ziGzR/52p48lGcIkSH6aGZI78GXEDqXFF97+
5goUPkFz1g48SV2iVRLLogo4jKUUGdLbxQWyQEr/qa/CB9/Dg6PCkdKjUlXOY+9t
7/Da/iYJ0BCnR8Fy1XL/SsygBSc6qglpdNRY4i01iDuVs6KH2S2NBZlhnJ4wB5L6
9qyGQNPoo1M5wezJELJSUV/ELtzzzvOF/h1GqgWbZLrWCbqwAKWVqo5nrHPuwiu0
N1BZ4M2ug/PczgKEY8dpujb7fOibHMJ/6f9ad9Yv453pp9benfX5wqn/5OYd2Mul
vbLTl/8AlLn7JkdaJEELk22L370gZPz+XAPddCyvOXhlIEVsSqKfj8pofDb6ELZf
wqdmz0aaydzshEwWsZYYmCU6D9KQD/T2EImwFufLaeYE0mDqqaCaqKeVKyU6eUpC
Zbb+8DyOyKJGB9G8DEfVHWeXzYS7dJxpMH5YgpnxPaGs8T3gC+/NNfqBvJavloqr
/DTw50I8YADbunOtiXmauZ/MjH/NmkfNt+qrl3ixAUkf8iZOzhduSzhcXvxc3VGh
jD/cmWaaoeQIhcdLU9Rk1q5ff5TAb+q8Xw4jfaS4pezje2nSJy66yMhl6yEDUj33
4P89idiBuL20tkoR5XLii7xH6mGKtt64v6gMZrJJHHTsC8SBnOo6RmATIAp0lpYG
qjekvnrnX59Iisix+YiANd9EmN+IDBO4tNhDB/2I2YsaQT2tAk9kvLT0aDkEmPi9
2NTa+/2peB39xPDSblA7FITHvXx6UhmTqQ9JdUH9BvbIY7iExEExZ8rJ9pvxeuQb
hsC3jXfmKV2Cu2TpfH7akbUJ3aHrVO9a83XApYCOTe6m4JGv4vr3UuR9jY7a+OwB
fQ4IKoWv6UjAPPCXX7WoiuyuXycATkfizDzvAuLWm3Y0F3KrtwopYDN04fyMIF6V
rGKuKUi6c3RN6Gs/qHYLTTu0SwHtMvOLltPg/XfmOO6bXoeeJQ6waZxQ+RKjmzy5
Wz5eqJ1aCTm5t01ySYhCQV3VkW85C2/1Ik5l7EG0uVUouzNrl+jlbpAH9HFu5q+o
v5AJDVnMGlqdX1F1F0R5/l7ASiuC/63XQxK4mjsnBWlEVAwnraOP4qyi71P2/14M
HWrqfCEV7EyrxHM32tPydwvk8D7YB7FMrhclgV5Ose81ou6L0nFqvJB6Av8ya5L3
eU1wwds3AwkGNpTxqnhqmkb2ABP6yDt7dbGWEZnzwS3qaTKAWq1Em5gejAE0CJGd
WTAiDmeuMkXSzhu1kzzeLLUZIwzzCiox3UES7hJYn9r6KeOSqs12nV2giwT/Hv0e
7Dnvc8g327RbmxHWEw+ANT7ry5M8wvbY/7da1xQ8AlAcLVcyYTyEwcz30uRysUsu
n3LC/kAU+KlEVbMZwajMykeOkfLTdWzPwMXRLPK9SZMC4wTFueZktJK9bVZoIpWT
aYqJxbWW4T4tEOWR+DrGwm9ejLmaxCQpXMWkuj1z1EO2TgOb+t62+D6M3ge2nNJv
+mVffgY1KbMxP0rO/OhYTNE6Q6JfNHVK6vGpPn+jGKt6iXnrkp4wD80AXtfN6/Is
u+DR0x7AXIUWy4uZ3yVhN2wqNTb6lm8xJ3hxILp4NbJKBBpsMhKJjj6Io+VDMfC2
Fg5Em8gIqvrM6o6KvmUWf3HIiU4YGibFtaPRGtE8pYh5BxwTcCwmNBL/WzVOqUgs
axB9hFuJCkSmvU0kFOSuOGMB91lp5A8PpkRGFMUT8LDZBIxwiNVxXQxy2u1ubt0V
3XjNLjNdHKMgzJ7AJ2Qc47bdIPHq+/w4J77WvnTQsx4Wly46n/uNwBOErMWMtYkz
oydqMQfOqFCGZrMUYTwwXcRsaV6fpHDI+aYnCZ69r3Ht4vv4tKHLoP5ulwECtuRH
4U852U9G1WxttZ6qC5J1c1VmWSmjWGP6yTzvzR5NdwNjF34af4ERL9Hu7hm8+Y4q
iEp8aNfoX5LbY0kf269ASR5p+GJNwaLd68CEBmA3b9dQNYREpd/zF0NtxOIRV4fB
BqRl6wN/LhIAfX7RgZpznkTiyoG5ZdOjTMoa1641+38sm3/CpRX/BmOixOLsgA71
fT7W1OEE/l0xN5sEQrQf3UEN7uwyNLrVVcF2JmehGq83AGw3OuImINbnwSeq0uqJ
NpydFKZa7osYwDTaBA7DoealMEfyoPjH1htVy1LNGzTxtjFGDQUv8rN+zqSw25ny
Kbw1ZdPN/mD/OBBwF8by3c/ozxLadrtBqOdRwajPWBU1gBGOvvFNZGH2AEfS8mJr
xBhhH5iOJogzEMg6S9ivm1qT73XLJeEEtfMfi5hwFZpgYPsBzkZBhuUV5pBNwFbZ
ASpAPQgco45iccyOI/owQOfVg1Rrvn62IlMVIzLiMon6Ngm1sRbI5cPtfgrTMbg3
y6Vphc9DmMPz2+qwf0Sv8VmLTyK3Xoj+xH4WDi0bWVcAq0alx+4vat8VbMVkJVLj
k8e7xR8yEmBfKP9s0tyUOyU8Ov2L+CFJ3/nOinbSnSf3K6Y+MZg8QGQJ7MfLazpO
YVGGMUJOO/3Z+zKvkY5v2F2jpdaJooaCCsXQLx/2YA4na4XGGmBh3cORPsyVpGz/
tU4pMh3evrcVbDvnPtmdp86Hv0gouGLQQRZ3q+BcXAARu7PbSVZ7blMZ2GfrCSeU
Txufq3bJ0MYTUQ9/EOj46PRdcz1ZfKZO0ZqFvaHP91MxWNpUqofqAvtTvwWJpFYC
QlfsrZJZAOTebgatH3uTpZOlUd1ahlCfd7kCQ6XiGlmwytZ6XYnYmknmjr/6Ye8Z
QBLA0kKqQ25cN4YvoAFasl7cqaAZwZYn9iZUyF0IKRrC2Ws3XBHAoZw4in0zgqrK
ogk+yCbsja8OYM5uqJc5wn4gCkAX6hm1vM067d0L1jEfeslS7e5hbFA46tpsR8He
/NAgNH/Ce1FmtMRsBwg+zTKUZKCFZKEB2e6qpKSh1AJv9B4npEIqx/6sqUzwiCBD
0ZMkZkSJRUqrQfgUJCRyXubjg86IDeJt2A9twTS64Usqur6CFRWVBp27xk49Q1ya
qvAxdDfKR1masqamhCuTDfy1zmAMCxTVMiYIqC45WGzIcfeWp483+dTa4AIwqGGP
7xXfurMDP2bYyC++91D7gO03XOXfyZhwnWKSqvDlgO4qj3o5ZHYzJw1pKl5zOu+6
kMN8x400nBSSDmgXKOjd2txKSOC+/nrAcUF4EB38hacNNhjJPNz7IikrAOYgJP29
tPCCA5TCj1IJxWdtzMPwo0nUCThLDM4qw36Jp8s/sYXMpz5DZNeJsAfVkSVwYKFn
bVARRVCrxP7JOb8ZyfHmy7GMv6zeCy81JrtBKChIyMl8pdXV8e6TiCG/eoetsrCG
1n2ibiChHGEuWSynoiuZ69c1W3YJD1WwrKxc2fE/30XGD/2Yr8R6KV3bj/aBzMa6
bqBtdZ62LgojU/W8qIwoqeRcSqnSpXT8/QvjWgRiolqhJITWN8ceMSxh6D2Os8r4
Szi/QQAfNcbofpZwTHiJ0LSw0AwV8yQVEUeA6Pu9WaLKVU9UlXW4HZgBkuV/JtwR
iJ8hKGYR6KO/uM/03JjyHn/MH8Dt1AAOnIZnpjwRa1S6iYv63gJiLfLrwGP/YtME
BVNmqn4asWdW7DPs2m459NOXQiH1QcVqNUWTPDLtQ/+POslJ9Oe+v2VvwT260aFo
4Y/r9dOGCEy2yLB7CxT59nBp05lSW1ujU2LYoilLrvsXhWo8GF/2zktcVB7UPTzy
//KBXKyXA1Ct7aZTRIjVW8VKF+Spa28kMsg3TGZ8TCGMSNiu67mpaFFkgP30XI7y
8iXugcmoBndSqu2Ke/uSZveE6VW8NnxTvzzbJW1eATrBD/1Vu4y5xgy9r7K51XX5
hyuj8oC+Ifgjk+EgVCKlpLxVX+A0V9AofYQXsBQ70Wlp4+mpsohabIFDE+qFMw2G
QGVtpLfDTZmKxxZBSeL0/pEh+gIugcfpr0fwnVkhOaN6tVUxO3Ze9JvZB5hG7ud4
X7gwglr9FK1MFAfIBzLnUHETSmItfJKHVfR4zwmnbypB/AP/ZZU7w8DVRTyukTHk
t6Y72cSrWAH3qifCgwG+GY4xfI5nY2vOkFB8lObAynE0q1j2Q8PihlcaAWegjNti
4TPHIU1iQ9dv92jxezxB/Wg2kRf1IUYeKEaWo4G0rdzYyEfbT3HHAhv97ijetF/b
xfLn9PonpVG/jSKmxNdIwFiZAQ1cH5qTB3lpFtZVdnkwT1eod9pJTR/SYRHWL8da
TebrRrRKV2q83CGHG0S/Q2679kU2Rnr/EgK49y7KzJ4IvV60EtRtzl9sZ6Oj6D+6
gHwJDcR6dyr6D/TDqv8lH+1x1mA+Jf1TjOBDqS38arCM3HOMR8SsYC5tsSxlLmNB
k+fCBaB/nZ0lw3Ji6jI3VET7jMaufQDPyW2DEQu7NoJx7n6T7O+nYZCnmJox1Eds
uAhKCSyhPG5z6ciUjvhzl/ss9NzGd0dFklr0MyEHd5/vxXgCETjxjZQdS0iwB1uQ
mJzG9C9DMudvXwM6y61D5DQcVhGyutezxJ2AEQfbFZnbZVAds4IWfT4q2nElDXp0
QcK14TWMaQHIC5aeFex0Vwi2P5/+CUXFZBhQlimOWyRewimqGARLG4QWyoS5UXvv
lk7UZDEHlvvuCNBA41l7MVFHb17pQsbrQkgdzE8VWTMAQEqzoHqxB4lPF3R79Mud
ToMUAhQd12VjXh1KOEcu8MwG6QJpLsfnQA3S9HanBOWdZZcZ1y2OLkCnWFx6ijmT
GYzW7RyW6s8fmSk7Aex9pLAitWbANzyxWNXNq0jMPqUe6imdZNAkOtwj7wwBCApr
VmyFzaI2OU1BQQYBvEa1MHw48zMxiz9ZmlVenJqv6Az3QFxaeo9BI/sOTADxmmfQ
IdaJm3sUyE2kJ0UsB+xrDQ6lRR8Py/A0XVacYeSIbnqZ6meDa0qo8eauaeNVXLDD
DRwdDYgGRouGkzHHdBxAuMknjuEDYhaCjzUxohDbPNBmxkT55Ib/dEQEURYvUsna
gfV9Q+Vi2Vho1I5i86TTLfMM8pzH/mjJioVpJpr5+ku5o5nbyN/JLHykLrWua3RB
O550tnXY6EjuK+AZNS0ylNcPuTPkegLjqP492ViQs1WVPgX+f3RZlioDAGyiUj7W
7BoBkgx3e/yG6/3wB2epoDhf/zZcUkXMkboxnXh8pJHw4sfEsnOporujKSn9CeJ2
rOFDkTAE6sHAk1XUZsobf/lmuzekf9CHi4SKZm5MZx1K/daTVNpxTBFzCEIweUsv
ixfeJlz3/Pt7eY4Ie5I7OvWe2C4kFmlZoNQh+gdGRC2RWrF8RpmigsqHajiIR7YC
HudLPeRYxSpMvBt9IDXcmEi0MvVKR/nl4WOF4YBMzDd7Q5XiVFYTyb8J32WQOSxl
ew1X14xUi3OESPzo7n/qHTSo5P+BqXoep1VY+32s1K6IamNJ27NULOLNcOswGGQ8
diPuTlryUHuC4+oaexlp+vmtj//qWomcVpDOTlIhTeEQAn6BIeDRkuIG7p/gBHxi
vypjM8p27h+KlczoNhu4zuJL/MenKfvmvSVPCVH24pdV8jPVwlGtiGn23KcwgYqB
d0QtSgi+B8iAiwbw87RBtX+PF6LGKca2x7HUeZB9aqnsspQc1wUHu6PpRPvllyLh
JBS4Ba5NQqXYg4MaDa1k10VKeytw5B5TdglGd/uWTWPCZl6iZbUXGktAaujCLBm2
ecM1kyebyNod/CWbKhqQoFLxE0WbAF6F1TKCoXFyNRT0zdpS+R8QdORbwWSyE9wO
8RFXgcm4xlks1SUr38rptd2uI+nKfwx56vexavIOFCVWMCX89Ummh9+Pd1pVYxuu
t07NDaZAhig3AmJJg1yBm23bkfSkrrO+Y4gAjQyNaGCJ+OioiW3+kLTfhhFp+po4
OtByhhKpasi21K92+9WjDAvGYHldvT00kubUhQwrB+V46rZ0NgdYqLYBCD4onHzW
rubj7giktKMaPQBW8OETXE265Tv1kVJms4oXLaUiWq7Z/f1Pz0EB7FqPgYy0fNf5
yjOtuDIvxOEoJu25cKf+P4aJyACGdc9OlpfBu4sq5wo8Kc8jcDnaF6K/32TKovA6
kV0s/6nHPsC6Yf4lf0jIsc4VHk1ik9asYOOy74EBoV+ucHu5yT8bU8RZCnvt5E6H
njYY/RBEHHeWYoOJVEW81FxabZGuELbEUKpjXZ5cxqJ0WA7Z01iHVQDe1uDAKNeA
ZFoslskXbIzBvpv8bofa4MEoEN7WKxU5k4yrWeqWcG5MDKsyDSlZmJvaZolEXmHH
GjIf5jB/qBM8PDiwejtcF7MBK/6fbuZZjdBs+o/a5U74SbOhHz9KcGRe4u4rENkm
bck52PZR+O0d4Z2atZVEbm0RGK1mlWXi+e/bRZDtDEmvo0rM/7CWkSFEAgwHILz3
VaWa0YaHwZG6/FgojBOO01aJTjOTs0Vmg7bN1V8EZ+vPSKsaVU//fWssJJxdAxsZ
CzpptCwpDCu0lZSWrsqpg9DHwWAiq0sqwNX7e6GASHzGNCK4jLJkNbAWfndgmt9g
zDWnGQnWhDJABNl79/ai3R1tsUEQRnCI23VjptCsLeei/tPlKxwd23yAu0rhW2ji
tHl1+rH3tu4zpgoSQifkOW/z95Kq7AAAecUqXnTc8y5+HDmjp3jRIGgGifFsniRJ
ULPCG119hJcqBsQtR31XSYcv9uIB7tEsBtKgSPe8Tkim2jxVbxwY6ZWlkmyfvVGy
gXk7VxMO05+OH7s8mwpK/ks7/LaOymKZAueOT3xP2d+p4ZJjJ380GCgouHobRpBc
XkhDPdTzPwvTs84kHVBfSK45p/88HyMdu/4JxZethk7kO71mRtf/WiNhcciz+OZv
I9dn5CVKTNl5xX3kX2aL1f2aZopUpCSyzXW8Pdo3/Prkg4ct7MvauDUmQqHYRd8x
9/f+t6qwDeFsNyOdKZtZwOzQjTdcbEPcc+QEwG4tdHTCbjG/Lu6Y33Th55phhnt8
jSiUQl01B2UfEXNbYjlhtG9uQ0WvWpQAJ8Wig0RzwglFLu2ksiFTcFn69d+F0NKp
gg2Td2vXa2rUhiVdr75UWf5v0FygQ9ZaoaaeEKhD9sDsODFuSPPnUiY3wBjNU7DH
lu/TK2E/cXYk1EpqNX01Nza0ojVD4AdlWIuJxhOosNGRkLrshYfTjOARUd7t+lEH
m4+SjA/WDbP0RcTJ3hYrPkobb8Lq7/O/higdVJxuaU1Qokbk3doSyUgMoh5u5x/3
PqFpmy41fhUFp0Qh4ANaJuBA2ynVro2uP1XhJrfDU77L4SOZ400L6BaEKqzdrRb1
xJJc4HzMC+Xd6ntj/qiFkyoxI0ERj5I7DNnMSvA9bRkveVDXHPc4hLx2qbFhzOyf
Xc06FNmb7/z+LC/3OkOqW6vpzOm57s0eQzsC6MfLttZTtK3YN/zCTcuQduDOUDLg
jMLNOyG7388Cu/MNAXAHzynuMwz6VhN0fko6IKLLbUg4KO10GmC07llUg0tr6mfV
zMaybDgx1qRi0mJLZeh7ByZkmhqpCDISLumMozjUAiCL4Na3kr02kZwgYwp7UqII
uyvXWpXhMzjRhh4bZEnQCBmgbF7pxwLTAkqiBfd1ups2nZnhRg+pqiC0OqKYX5+W
oVfi1MyhemKtCKNVs81OwzTBGEcLyp1Ww3kwcasG9Zq3zvg3V7v+cvv1k0SOu53d
zx+D9XhWDQfR0KyCPnfw4/Eju0Cl2udawQ7PetNys49NBCXMQt1vt2J7mRNcobim
6FzzX0BoOYX41DRYcB2Nw42fNti3JAzWdcQS4f2ksIer2D4tRPIHfOHdAHy3jvFo
nQ16pUuxgQd2vAGXjcZXJ4dIqiQ+cOlgWKblUfiP1nfxzisnJX4p5k2dtBmmeR9e
f4fnflGQIN23wRHocXNJg4lyVICam2qpk1WqBEhFeQ41t9KTjSnpDQvy+xzzmlH6
8P6vh+NcESC1dF0eUSfxHe4Znuuwf5YEU7P5p77oMCEuQjbNV3w6t7I05RR6uFVF
4C/Em7w9zw7vJzRqjQF6hbq6ddNdHthZ+0CS8ouhsyMiJgvTd6KsN4rLoIK77HFk
dpmflblSZPV814rWUvgvj8Xj94LJqaBbDaSWQ/CFAEP6larcs6SLvRoJp4zq0FQT
3Ztf3FfyEE+TEx9nGb3fIPMO0IVB/kH3pUbYknnF2I4+S1aMfI4TMDsTG6j4LuqC
OEjnOgotVendvIR4ES5d/YydKJDDqXxGO0NStc+4DVXY5Iu4fkQla5jXaD6oYhFG
oKg54XaS9Y1TQ/zjotuIzQ0pE/rm/RkDz61J2iK8MnI5hFK3N05GEbQtIqd6gOLy
NVmU4o/seDjs+QVRsbjL79/6HMCiBGdD+5ZjzD+jZ8luIL/6n60tvdnl3V9Nxhh6
ILtMY6HABDwy+3BtaCEcBlhuD3y5vx+82Mzaj0BwxvjzqSGONG+uB6rLmC2hyIns
0siYROCMAQEGrDZ/wZeK87J60hk+9x4/EEgEFr3hBt4pkT1tQd16X55shMIZrsKD
QTX/MO61GMFVUIF+U/4wdf+JYTzqeWsxUJkkUMnqKBVmPsG1lqc/8y3WlhUk4ZYe
Xf8THVREx51G7JhCoeacixAnk5SHRpdadVXHoDj6TGh7yPmPOnRwpY+wQhfAZntl
QWE7HaGHy0TVYRxzcmwuznR6Iv66CEjP1fEmcaVRmNCqLA/rT7KDvZ4DZcG6wsh3
xpSC9P0rGvsn9JxBrz5Csk3vx4MSEupYW/9gmK1chCPyKWNblQ4nJEYgKw3LZb6n
seAXR7nlTiNX0cZm8QESOLPNKKwARs0ETo2tcgS46tqOpnPKY0+inm5T3cUl4IrT
2GrEtX3ZhmjYfSyBYKUGhzAgG5j8FE93NSIEIFiT/0j1rBzcBebbF1P53Aat3VCp
p7hw8DQlYalWO/ur9ZL3rJogEvJLSWts+hKBQ0sd0P6MK5IZAzJfWPv/Kfs6wMxI
5cwohP1g53AOOmuieoGx9a52Tzc+wAHmxQXu2AUYNrWzUDoCPGWdHuMbJT3FjBeD
FmSQcVsjky8NgoUbT1UgULcZHcGYApQgkMqbsSt4sr0VSsbdZouTc208EbVnrKK1
taQKMKsJrVwE8z+kbqy+JxKgKHfzlBbMsbQPxw6HDkdwt5/n8Xj7bUpPeLTYP8K2
VSUALe7uBJZ1VAC/2JvMfWiVgt/2UfPbVEpYRrsbQFsCGl/nqCyJLGzG8zICy5SV
jiho/JWDPKL7WjuZU4SPuTHYdZOBSm6gCTbKV9NkEdS0Uq0IeiBvTEfKTau9VvEF
aDUPbuEYxHG0YBOsItgFEZz+BZNQft0tPeFSuySdeb7VpaHS5x48CcpLvzlsGxqP
sxagPK4MQZxRKB3AxIM0aBMXRSNvIZaZbusZz6Qs5qS/rFciSWNDdJ8VWmoDguo5
isBDhQkmgpGMf0DuwM8DkvlsVJXYqoPNaYTrU8QiMNzwxyn86MbJtjq9DOpALPgU
LMz2+PsvHAZKdAjOc8UlDoPyYfd8wYI44rDMyFqoSjbTZrCsvG81FK9mKA4nJgwl
QPUjWi2ay/Ra6032Ae1Ime5kIZ3QZs5xKTAqH+PRhSZNhnUTJnkBx4gjxzOiBnNv
7YP/FDrlG9CBXWJA38Gc+li8PWrTPC3mnzFzLi7Ve/NfkNvMSWQJvmuRCX2sQePD
6gN4bbIPI4a7ts06o4Pvf+GogQ2Vi8xbGdWQGfsk43lTrGtFe3MRBBlkO3CoPy1I
5EbCFMRP81FXLizTufkd7KeCSJBv6LS1ss8Hl2h9w6ppoZrXIqIWONT4GvKCYfmI
Iu4dCkjmUQUI0cTdPjoiQ26XdRFuPGCk/jl1PSPRtCy2NxTXXQZI/6ZP2ofyjFN7
3s0AylxxI3EdpJZBLapERE77CRK8tqyDnGFIdSobzLHqWE0ekOB8UdYOF2Qnlhvo
AAQF8d+yYqGEL4RZ18dCF/nsepiJPJ504EsEpZIrvFCAHk0jT/LQxeMmYr3rECiS
5DNsr8kbv0oB9Wp8d8L/zyQ1qekbLkRw9/z6SN0tdAlqfP4MnCBFSCQHA1whAzLP
lXq8mQBgcwN23bVpnwc3iJ4fmsXrIuS/GzbMToFf+Gk1PjaEb0UqS6tOQ9VDfU2l
HkCh724MOakZSZDlM7BsRPRCMtV2h1fbNvCof/ShwKA8N7am5UuMYmVWDgTgAvGh
QSpNnA8XvGuLlfD+90opI1UrP5cqu2iU3l8ZLOXpxBifXkOd0O2cjjUYctYp1vrp
alRNTiyFzMWWnRy03l8q98BLKB/OBLOfTBzkm6mY7eYVL5BrzHuGOUMmznGC8b8F
E/dxX4Wdk53fd4pCWh3q3wceWyb16A2CYTtTD3L5+dRirjYi7aIFcsjwN0REFGdv
wIIjSYldPTao3orZJRqPJwu3WbFRvsJ5bROwS/pvQAIGBWMB1HUgy5xJUYwcMWvh
MNfcY/b9xxz159sCKU/NS55d+oNXIrrk4CnVysKzt2DZxhPztK52tg9UO+2joTWB
G6yQxmdfM0EozwMiUx4U6HxosryQW+ANPD2Tw7CF2giTx/hIlYvyYSJ/5Jb+TgP/
kdSrvg2dEd/hXyziGSusbh/UgWYxxP1DJBYQiEnwDw7lYNK6x9Dvp2gdZpqZcNJg
Bbi/gx8mpSpGIBDwF0BlgUGZCh48FdlA+V0yauRY8+DSnOQrJq9+ebKF0ti+sk9U
KGEmzuSBxls6eTh4T76sv7ZWi34+NRXw+uqKJK0j0Jwk/GCHQJVZvcswZRDWRP76
uQn2UGlc8QyTvkmgYW3Lm3q68KrK9v24qg4H3uJpxdmRJcD0KNihPSxzAaww59+2
WfFqV/ylB19DfZSKnK8jkDnafE6ht2NlaH5yAdBjcgv+gDsQwZXA5Fq1vQp39fPA
HTeUTt8OpECgmmteBm4ArBzYbQ1/44dQmc+nuyXyUnJh27QV0MdmDWwpi6fAFF87
sFVF3AZQd1uqGO4jlwSYPwqpMgnHn0vkJL3hYyHw7e2YD4NWZexPR/STS0QnQwXX
wPnhhWFN0rQPYYgx3ioaR8j31fTGKG9qDYqRHm9MDke390YAQ/s2CuEr5xLqvJfM
Yj1qLPBHspFJQS8HPGRD9bb4u7FTTvkNqh6jotHenHKPHd/qpSdBs4SdSkgO2Wx2
SmQ60dEs17wj8BW+/tHsT4X5j0Cz7gIrhYZXyxRVT14+3qvXGPtY04MYPJeV2w/Z
e/npN2uXrm3Pf7VTzGChZyNEOtGMMoWLBUCp02OtAA2hlY1INpxcO6T7qjjEwy6j
vIG88lxSayiWj2WgJdY+1nWI12xm0T1VedeHJ/Jyq1w/UOr7KDjVbDimaiTnwwQ8
kpobXb3ml5gUhcHugiY6lOjgG9ox291DYhjGhL8VnniJfmH3jT0d6t0hErYSLsil
6zDMwQxXCtZcQWQxB3h8bPtwBxrwSOzHg8CsR99Fp9qLXqBlAaMRxZ60nwpF+ETN
KPrxk1pxzi/bbOLGAdRqDZk4C3xoxOSSrrsp+eQ1cZF6eXvF/tQhB0GrYP6ylWRE
rF3oxAP5PfipPOksV0TR1tNiPP5eeF/7C9+qL7nMiLzkRgOVRe6uzyFmP7tL39Cs
sFSwccEXMVmSLCevntJVrF9HcwINoB0GOcqbRalb8PWyPwuok0jgjPG78/qaPlDR
Qlq8az7h70R1fPKKLh1HJOegjpoSpjoS3UivB8jHFbIDK6j5MwN0mLSQRdRhuS2b
bsH2XHEF/3oANoUOaYI0zWwln4sGI6n20m7SpeyxKZLrv+JqQpsIYtnfD9P9FFFV
FZcH1Rsb+2Rel4hq1FxQl5rGVIVyQycjxulrxSz+u9igycW75M+2eyfFz2PyTbSa
q2e7JDLg1f6W8SCbEzNlgbo9IpZNJ7yxCbuXNCuP6vRQSjgn454VC7pB++cV6VyO
bfIiiwQTh9H8MRRtH90uQg618zTZvE5e7j1dG4/zUL4I6ow/LINBrYnqeNDKaKRT
3PD60gitEmiHjBuBTHGLwuNOu/hccpicSycrTttIenjx7/l07uEqpfFsR2OznwV1
Or+ESfaBNaXCvj1HLIyX9oM7Iw4aewG7ONePe/sulitGdPSpduznnNX5WoJxUCkj
vuOWXrSe3Pqgpz1tn25X0tsiFycpUiyO0pwjRnkdy1tTTZYeyzp9+3v3Y7j0M4yZ
clcXXVgnf56UQmMSx2GnyXWc2hIRdoAb33HhJY34gVjVAlBZMFMis2zYC/zKYMOH
/fhfp/ofUrzlKACRqg2S5BLL9SZ7YILjQj2qPrtH3+qa/RfxUf+1gC6w+OoZDcYr
jjGpbKIRuQs8C8eATzwGclkgOZqTxgcnr6644nG8iuwXXVS0FnRNOvi0wA+AfriE
Eb6w7V+rAY5hTXnf5wqx6eY0nP3idbW9siGj3NpCND2hNk450lAGRaU5oN8YbaRX
7OGBwTmppFBgQ4NikSe6didvlwEXHFpoU3DZK/CUjEa2iha/kJVMSOvtENKUf4vt
Q1FckXyY0/HAIGPmciRDMOsWAqf6BxLas89ydeUuf3BUnyyEQQX96sDa5QzcuQMk
EhaJolM75FSZcOFWAD16yGgJnQzsGowBKkiznqnpNYEi37SjfgsiWHZ9rzOE2QmK
U1r41ZG1LLTvBPoeVaushffYImj38owSP2wQN+iRYkISr56UYilNYp3nEmR8KMw0
EwhiVQsv6nQC/6vN47SCXsP5558R0YPs8N83sMWJM07TgHzfecmJW01Xs5FZ3wVb
S+6P8sQ/T8fOmdtRITtsBEZ7AIXFMxaXIduJ9BzQLlYhtYdgOpn7m3TnB0E7PMQo
ImTiB3G0HSiEyfdJqMaS73mLE+EEFmozbpbQx8DS5UZ53qpH5rf+ZwRxZ0zonT/1
QHmmyjg8r5upB8UxRuLp/4oRcIbGQcceR4C8KA9gWwL7nVKmtz6DNwOyvQRk8WvI
7yfNvBQAanoT02WNTXfdOTldo7ZuNz63x2RhynjRcT0L+hM1rwyvMV8l7UyISukf
NmUe77IiBfziBAi14xGoug5hTneCwxW6DNvCqk4WJTpjP45yWCQ8E/BSXBgpgl4q
RFLjPr3BHy8aBaBp49oy0VtE2ilPqnYK2S7Jwco7+PDLXLXyFWoVcq+YZHKwMxOZ
IPP2UAkUgaSGLxT8JG50oQN26lDxH32erMuAa2RPmg+0Ha4/rkyx8GltET97nef8
0TT3+ydKw1dnHGDhfaucrrcC+A7sYlM57mn1UaLS5hcfZ4eCgQsnJAawe/5ydt/A
ibhGKsaJ7JQFquBJdxxSJWmWxbbPPDufgA4Vrfh+ZpCUvM+8/a6gyir6g60zVBk0
SJoU5iGVEVC5k9TOWfBhELVuzWKd/7bhVnQlX6ObnDD6jtdI1gOqsTpy4f8ZHQtp
St9PSQySEQA9nwRjZwCa8j+ruQIjRr3i/mdlc0FxFdbi+QvHCF2J/bh1PejVv7C8
vpCej/HZxh1vaRtkPlKL6F3oBoC7Ygag9RUc6Y9NHODRcA1VwhQZlqRJDKIoafik
UoGn7AhfD2Wn+uamsDtw71bM694XWjf4e/uZ21sF5vWPwGUXGfEYEFG/p5uJ+cl1
KEqEUm/glzg8pSkgyyFrdiyTd8yJ0C7+Xq69t66xQIFrmFEpA1QJj/p/szGDunzM
IXkOys1eb1yEIFv694Ilt4cp9lAnruzUFvQm4vqDIBtiC0ZtoQ9xsWX7ZRwbjKBB
jJ962ptpdbFaWtQkFAcqGQF8W+KCO77/GoIPColUEO51nRFZ5yWYPMq5h7HPzkGz
ho5GI2vttBFcX3VxzzOLu5pcwHzdG6QHBeIcQe65KLh6oPgKBJVgYwEru1rGZYDK
06P5bWnrH1PfUxr+2rE2ZYOjNvGTq/ysck3C7lXTmern18YSFrM9r3K30U+tNPTH
2/J4AkQO8mMDRmbbY9fByzjPHFxnKoEtxdA7mmGt5ASe2iz72hnyXDlNFxpCwrOu
f6Mm4jZrqB5CvnfIV7FCTW2ULoSjuxPnE+RTC5A30f2c/lEobxN+WrvCLQbYSjls
aFJUCP9Pl2xnb90xwdyV0Dm+BtWVjJ9vGU+6lEJ0x91Xqql3XjxhGpOdWEwpulUq
jTsQdKT/jV9xq6gMofDSr90cOBTovZhf7CI2wm3xQ1JCPVgo+ZThT1NIkqCSxz/N
rtEPgj4XpXlSxTg3N4c/eszoyhlhVNUUW2KD7bVYPpWdSWyOPdJFFDsyT04mVklx
YiVMAdBkMKOMw72LyTfLO9JnfIHWnTjDwD+3fOFWs+yFRvjGaxfGciTKsm92qKyQ
0vBTgaFGU5YOnpyRutn9rBMndph1DXV1ME0iJICq17FGXGYrdKLPBc42zl4KnF5M
pky/z9RoiRSpwxsqrbfWaNwcZuevltJzE9KilqKuaJs0UR/qlPq9jjwpj7XCxye1
kjy0zL6+8Bc2V1n/7u1P5bWxHHTFkWBEOPgJbBxxu+BfZKo+GarVA7zexy6i11oe
YG69hWYx6i3Pf6rWi33yBjgEbID4ionCmTNh/B8piN4Ewfr1S/INO740jCaG6Qb9
sfTl71ry9C2D2FVzh4vuSYoRaywr+RiiyVqx6yvQoNaswy2XgbZUjycHJxbIcviJ
itMvx5qIdLtESWcVxWp00GlO9pbzUG7DFhqe3sDpcwurm02UyACpexS5BR7D9jqa
bsxTWggafuHUORQysLvHqf8HFwqRL2Dt07w4XR5huByp2ODjGzaUd6UHnJRhg0Nl
0AGr8wg1sU8D0yD5PLn6oPkP5Ehmtyxi/euU5/2ThXyrdyyiRQ+PbyC7RWX1iqSH
ygUoJWVues12aw1Ox6PxS1IjxPDOiwXpnHURPryryIBmPgpz1ghUa+/iDwoh7FKM
FMH8B9dJm4nB+OFv9bCb5I+1NriVSQ/p/iS9YoGl2JFymgxyIAW66CKLJF4YdQtQ
74qhSTQul+2jHvW6eA1bSt6pi/Sds/R4fTkGVKgJiGRV65izYF3lxnxP/87aYaab
c+EdbZGgJ0IDFSO1kitgg7yI+2mDuh6bit0NiJZycIE5Id4rruaknO4LhwbhiQLz
QJB20uWCLUa+IcL2Yadsar5I0rPOIZgZXEIfTIGLegW9bZAMtFjOn33nQPE6Gag+
7KMjclsxiPvSjqJGe1x68sdNvSrvNcxvcN4umlip4jfE83dXoI+naX0HIkz8KcSo
csOBhIrdgTL1HrCajg0sdZrRslGR6nkejUJAFmNG+aLOCSGPFcahZrKfvIi1sgXM
EgH80cinyX9xSTRlS4VkKOBHTAUASB5IGFOBS8YlWHc5J181KE7D2NfxtP73yQi+
yqzJfSD4fwiVYJxUm8GRXp+2osRBSLyaKjVXzcLKw23LtW1ZYB1QEV86nlJuobIK
dxeLdui4JXWjko7O05xY1/zdHkJ5VYB/GIq1Xs3Ne25B4nvWEu9BrjVvbZgljWpI
vjKq+H/LpedbYzcKF0QT0WuctRm7269CCqXNw7kCUsyAyVOORW+m82EqHkSRB3UZ
OvybmmTAQy0lx+kwIAe+xYROaOir6ZPGjyvG6fZ0C1BUuC+FQtnMQlqj+KOCbAX2
Mk0AtClBiH3ulcxl1cMYmfVJzLntXz5oBKGAhO+8aXYRI6txigye1Lb7MN0ZHwVS
oOUP680IZ65zECnAoghmW9+CpDnPbVhne3+klgJ3pvrm9wq5HKiQbi9Nk72C6plu
fYcxHuCzgulN3+y+BN/MJ9Q0GfDcpxh7NlXpCFgPGfur69+4o8SMPeHAmOVpHhlO
DQLcipew/PhG3ETA7kjBkycHJB58nvLDxp24ZYTJ3yDFndtuxgHt+4kDK2WGFL9c
Lw89ORSw/icCiTjjF2blO7Cbo/Bnnucax/l6uHLNHQedthvLFu+o+Vg802BfQ+Ir
+ZK5m5wWyh3BQlHKqXJhzKObYizzWv1bm3f7y09HYvMemBb1LhJ3229FR07nJAHs
zizFiETL0AOgMs+0rnqbvHWDYwn9UwM87z3umn3K3tRUMpkoBgv34sB9ICrlNFL1
wk7bzPV44WLWI+KtFyiLUPnhNp1qjZdeehf+uldVmEphq5G1fGaZzWdMOwzXw7CO
WZQvoIH1OZzCdzP9iMvbnkpJq5DQ6n83TpcqMhNFqw6ElbvFnjUI7l7xBMh6GCtM
EMNUAc+ir+c0yovSkdgseQiE4l77lawBHIZ43TxeShluBZRQSpc8vigv8FF8k+Tq
+76R9INzFV+q+8ZzHRwGvC+cibKP9pkkd8GHbBOd81eN365kpcFc2k6gTkPRgXMM
YIjaoiYG1dm3pNLEqsW+RsMLUxvwOtGR1hmWf7IYylhQ6Wd1s5I4WT2CPXLtYOq3
vmRQOpOzdGdrCwVva4VND1EC8phrOVwDOEHMXEEzsvsUOYgyRFzg3R+9fp/u2/gK
PxwiuOl1zOMFGMtdsOwLQuQWszidSdmQvtI/S2at9lNdfmqFpMg3StyEmdijb5++
Z5D8rXvZfUwJPdY3dlQA7UO8h37qSAOoEcqrYa6JLio0ijwb8Z0+7ntBt4TtnIRt
PevyEMAD0ccGYQj1PHaOPKzcV1XqU1k0JPUwUKzZ4uKSojBCH74FPzrMvE9nZgnk
MCtKGFOm0rHPjtFApNz+y85RPQOnLxNvTYocgRbccYKZyMfiWo55D/RLTRchJdC+
X+zpyQTUX7MAmTdRN0w7zSpGFTp9XXg5l0JzleqXKbSdqJD4zcdtQP+9LF2TW30y
SxSs7v43URohHxHHjm3MJT8PBxE2H9GIbuBXsV5X1fNKBMnW6sZo5BuWk+jMYo7m
wxg7TRREvjZ46bZzrLeUviByEXfsVuIpK2fE6sR0wXoK1/86qJENYDKV2FyTRu8L
2aT+uRjruoVZN+FADQLisxCEX8KBJWhU7A/H6dX8m1AXhlLPJhgWE/dmFpTCaLpx
9fPqoLJWPsh0Kztw13PkOH+TZZVcF06cqqXsHrC/kA1aukp60DrRBtgTB+Fk1rFD
ZpRXDAq20gyKPJnmaSgxChB3LtRU6HMCKuILQLB4rhtSyd+WyumkqvqsQG9vXS+i
OK3vHc9vAtTGTuXbWcEg3KKHbSXZUDfXuGWWrYE0apa7rMJM6RrioT0yDtQI0820
gs8WqPZhegY9RL4Z+3PDG6TId/Nx8gIoPhG7t+QmMDGyqYmIPBkiymFwkI6QkslG
1tiaVHFMDRAkQcwqQNS5qdb/K6RaM6MToHt6enMjpgEYk2hSmZNhUocu65uXybaW
3LRJQt/8Z8KbBrJsb0SlMFhoQEmGeLs5/bKf0YsQjI9ti/8UzHST2QAkdC1F6+FC
r4KOq4cu9LFkHLl0qr45m34Bqoo3sZiAaWZN0Apv1t9e9d7JRJ2K/zOpIu7iMrp+
jE6kFhlE/hkwD2j0GPgC7zTfsYYpvaHZkCbhBSBm0e9iu9eHxpnajfNs4XQfKEs0
w2wzukZvHp6nbMSf2qGRgUorAx0HuZ+A+MxhPGnahIr8XoezkUY6kHLV5uNSr4Bw
7vtu+OtxftplNPAdyM/bBt7E95Bx5JiHepTMldeVWBjFXkDFQ3jJvWNx+V/GIRpv
ewSUQ5tbCFDYX4stuWEWhFbZn6C9PXCVUO5csZEsSm7YPVlTqUIfvH3waU7WtCXs
a/RV+3J6LaYP21BkWS0TrRhpEyC7paKJwjWH5Um0L+r5j7uxNqXMW32MpiM0FPHz
8bO4sxEPiLCP31ptEu74X0Xm+zRcycHMDhiWHUaJ/OkUOeol0qqU7zn4n9Q2S48j
ev4Q4vFQ35Ek06RSkkt8ShoPW/4CUbsv7tFe1f7XflgxOvMd5599j5IJ4/L/y/c0
aXZH44/AgLtiQU2gHhO4LCENoJt3pClgaPb0dyjWAI/9xqX/RMtVAmF8F+AqxKIH
85UpwDeF6i2kIRLI73A2xkNON4qvYh7R5O1sgExu/yls7p1zs7ar/Ygw0AoQSvST
vsoUmrAz9VjqIbkTinwv+EQf/5IeaMmaS15JYxRaVrFU66hBIOaIH4ZsQQbhz9fH
M3iXikk6g6RRxmD+6F+MEWiIHmBsEd+RnDX7GAO7oA3m5reUl0RY3hlt0ncGqk2L
6wbPwJvf6jRmcIgjbsft8EMUpRWtYtjwbELAfV71Kl7dhOq84oecKpojSsujg+zj
SkT/tR0tWz7UkN9+5He/ekHeFNkLPP3SOyA8MQCcy6d03i/lHP7VGBQ41p5bSda/
iumg69nguIGXBLGrlxLgq82DYbWKM7kp8DC/hZz4Xo2gog1z+x1yCbJoc6tApczU
oRKcq+0aovnXzYXJ+QgHEN+qlrXG0fwU08IbqsRz7QHARw88yRdDTeqEgO9Sx+hj
F86/vR5y67Q4Buywd+GYtGHcixOezrYG3evfELpYEFzZNB0vLQalbenuw/rtG4ls
Hl+0cR2tsvAe4KNIiNht0+vi1yHA9ViMCrIcj/QvAPLwTtkIMq7PQo5yTPYxQwsX
5K+n1/XLvSfg13hkdU3qX7Ryqss2lSwVfx/JcYBRotiBQQ2M4uqNK2ahFBtFhRqL
WCTxZYY741KnYgwrlcwOvaVUfSVI1nrA6CXUFKbsDkMdviv3XYrd1/X2vfzx6c/W
N8zVXdbMzdkhkpzBAZJqs/9JBPcin6xA9A3YCSLuz4EC0bQbQRAmpRTGfQvehxar
zWEHr3puB1AUvXBohaWLrf6DlvJ5cI/0KhcfMfjMbjmhbUih9UOADDWM+qOEmwKy
ftAUHJT4kWBZAi/F9Wm9T6L6uRjgALXb6GUAHBqkRCJH/96PaeqTq+Hll1yb1xAB
wNA26uquBfwZ2oQ7gm4BN7kWAGo0mMPZ0rsMB9hnBp228h/K+VxECiTgwl4kJWmZ
aXySOpU98+CqsVGtdncxHh+5j48jK4qZdfiTkNsQMhmrywcyJ3kmKwF22pSp48B1
7qhxbkt33JeHw6eTTQw5loKpQurbdyM7xme2XBokZ40sjYAcEgD2cM8D2zNwQwTy
fI/wasbEHwRTYGuEZueQtC32CPcx5bYjoluTViru7QGd6xvCpCKeIgjDEgPB+5PZ
QZ3XcaqkXQ7qUFgowxryrr6gqWwM9E9nQSkifs49sxTkbdOfRHmqQjMD5SDcnBE5
pHnPVDKWsUE8xSQppBMn/Rz3fhz1aNo8SInlH6klGCSpnVNSw5GoLq4oKd1k7h08
xBysVzKHuifdh4HIQOZoqpQKJJeWqr5wY0pUOc4TEpR+xE9cwlk9nOWKTI0pWCOk
PEz0/XYAgvzSXeB3D+Fv+GyyaAiaXV5LF4UrjZ+t0s/Sw1vgIcdIvX+DLDNuDCuI
eZT5/mJuFSDeU8y4UcM7dTWRtr1FRBqAhtKP6PbGcqM98obmAMUEAwdREuFoCuUR
rlNMxz/XLCiO5C8uHFpPEspDhfhS0Xw6mJFFu2EkN62WD0IGdrcVsErPMGH7kBV4
3S+7OeIqlGQ31B5qw+SN65Yis36MdayYI3ACj7ZZNn9D7on5S8GEBR9Dhp0PkRJr
X04ysHZ424uP5wxavi6NWvQDnKTwliarq7Nnm5bgMvfAiSWaXOBRY6dkj0KgIQst
J+JtJHhqdv0iiAucNQVWcl54+L3ryrgzVXp4mxf9jd5KEWEYqCjG0WqVzFPZeYCz
WQj0oxFbxDannlwdHhd2qp1vJjeOjvLYtYpU6Zld0CWnUV6Ds1fzv+YLU0XUGL+z
3RLb0VcTKsmbWIGseSq7p4JIvhBfaxhg3WwbTuIlrN4dBDUHtjjnOU2xDehrm+H9
as73ZMmYhXl7vOhQFrA4M8D5bJLwrC2polrGfQ6JyZSLo9+nNdhn8zBRTIUysBoY
vfAxVQTp5NSzkkpOYZtd1Xft1ntSzDx8mfwnGcLUtinMXU9hLgI1EkSikY+zqmEd
y0aD2NX+9w6Ym4xjTyVql/789jGVCeI+MZ++azmJDngCRSOey2XhEXGOI7I7m2Ap
QfsgXeLW79yg04joZjaR1cOKHd3+2CLqqWr4JCk/WZZxEB+NZqEpbp1lf0+sFJVM
J68C06v8fIayq6jeneuJ8KcUJ/7QK5I8+IdDx/EHWlAPfjn+hR+OgMPLHM1vdMPu
q6JyLkEX7JJv5qorA8B3/8zBoQ7kuKgND4LjD7PYgT+eBMOo7Atz+PSylWjpje/f
xbmsw/NzMk3GD5x/TiC+sq5k049gdmCyPIEo5vQvgLocsgL5qsINZf93jNuFLxD6
G+NcNIHs/H3VlrOegNBiLw6B9I9ZsgqXEannBQKwA7hJ9B+nN+ZxcfLt2rK+yMQL
dkkWHlD8wdSivJI5UZ4nTXVGQuQs1sSG36/iPJf2xBvO6KgO7IApu1f6yubB4Xp+
RmOhPeU7WoIaIqo28CCi/iLy44uiwPLheoZhR8X8cFZyEUHPGWjCqmqC7o0tVSDp
5YT+OiGFtIO5oHVr/ZGafM27MNB9Zn2G9qKcqWwM3uHIBNZTxc4xIACQZwEr8VAp
rv5TRRzh3Cpl72cAilXEGhhZZMTQdQeIXqCl8+OAgxa3nR+fXQg8a9l/sQEhLhdp
f9EEB3VrFaS87uxvlOzEwaIoDH6f+ks6q1rDxu3CCJlaA/5I3OqNOXOOBSq2Mzqh
jQf1DhQki6IacRht8PYUsBS4MTS7mNitDMgyEFRGrFyiyzk2kPyto0Y/mfZx23ad
U7AHQK+sDzvHarhc/OUWhLzxNfvuPjYfmx3qSNM3gSOqMHy4BsoHQ6WQF+33mxVB
IVF7HMvYiHglyNsfYkfT/PHx6bjCzd4Xfa4kAaGH4i/IYZn7VCiBRtLuHuA43YRL
f+iXxDIn+Dzo2dotc6f80R8M3fg+gOQzkIm9eqAXGOtFPO62H6RRCKlXuHnNnLn0
7e/i0XGwUwIzFb3rOdsdJFS1aOMI3PD2zGl9HstQjp7XwvUXkIHgx2syMxzKETmq
DJj0cskoXYn+1h9kPhznDhxIBV53UIwhmNiEDbsPiQAsZhoHOhlE7NnAQSFu10qk
x2mztD8Z8p44M+yiJcPbQZ0QgE9VEYCBt+Ls49T0ZiAYRVLzBayh77EKzNiyWbbF
6oC8iXLuiQLdy8dHWd6MD+xGqDLNdFV3+iP8NzUD1MHN4mKNILfLd3GFmRQo8j8i
1N1lYwYJ1qaam8I0hlWVl5MNi2FDmTAdkNxb3QBCIeeqUVTrJzStB1B9AaoO6xq2
6rC3fY8DPH/++Jxrj1TtKo0q0Pu2OZpY56kBi2WGxk8ahRZe4xB6AQNgLEHc+iZK
h8BfDlc5Nezfx7Xc+NKGd02fNeFNpE/NF2F2pgaL/uf1lM+3ivfhomVl0ptN+MQB
NlF4a/yclPDnb2zmD8N+AytSwqwqvUZGQdR6Ln6QvwuGR+A3W6mkdmhRaQyBDkSh
pXK0Uk+ffV6LdWRdQFs8CQ/H6zKfYl+Q6FsMVvHf/+6GYA3k8WS/ObohDEH23xrp
XWS3W+7W0gdGKtkshjpssxENRNAxgGAa6utCMZq1Hkxzu0TXA3QjvxieL1XTIoGZ
j4SnxAEzyDzcjJ9OR2Qz542QbnT4YdwVT4IPC4COXIA4Mm+LIylTIoaQAQBdjJ/F
OeXiHga99lGc7E+dkQaJdr6DAj9+OFQAepFzSLzdNTiHLDzle8NOLxI5WecMTtcY
Ds7q9/p/bANepvBCJ/Un6XkK2ppjzmXRGrE4Ud7ue1F5VT+kXBtunYvWTCFkuRgQ
94iDT5Bs+Q9DNUsKpNTj61GOp140e7deonE1Peu7jgZsd9erekECZAeclgKwjPhr
FIDhesFc4VfxYyuW2LdQOPrlZaJZTe4FV+mXlgoKYIhqTpsgxvmfxf1lb62riwCK
Nv7IDmcJMBXDhhX+50GclnwYlqlZPDgRUImdHjkP7AKUOCiMTkCMIjLbG2ypfykO
k9a4Zg3XyyneITlBqNdgUJXUffIDiZOogpWD8WZT0DPHjTMh7xnq8zueTc1xD2yq
0/yn9byVaF3G9HqWPGXaLsNw+gNBP2VQcv2qTXom6yGyDVf7MFMN5wBWGAIfNWgl
b2qRRr+wH25ORa+EcmrDYCpmyw+Y7jhSoGyGaceVrepLe0jFXr7p994WVPZ82EM0
GDOBAG2PZ3HLVZRwTtawXl+kMXsD5yUmj+mKKPGC5ZAAPOXf8MLc629Js9NCVuyf
EjXr7Hi3YmnFn3duuXdR7I87gioNI2DolysTVamH3GL8r+5+70o1syIEj+Mf+tmJ
qCfY7upzlKrZZNY9xS0RZe3SPRYlYNZ7jKfK/RJitVnpfptkkIKF74YfVA4OGGuT
LKntWnoSpf7SO8MwVnI+8z6T6lvns+FhB1TsuL1sPV5I3f8mZ3rYLTXhgXlOuORq
hwofO8lQNet2b+GrdGLmTNTQQmEYLttpFuHDPPJbwicVxnO9SBU+uFI+IBw1Bcin
eNevtkHxTn9fu+L9EaXbD32yP27MEnRjnoL6eYCfJkl7e/E1mGxTqKN1Zv9dSMB2
UJ4sc/qJlN2x9mbxHPFLPwO8GCpLBdzPPE2YcZo/k+dzu4QqIZLFEeOgaVOOyxXw
jgM/hTzqHgihi802r3BdKsFIg7CA9vGdAX6OhkLH4/uGCwlteeySKNXCxFRo5mbv
mR4pEPpL5Q4wg02jffFkgAFOLn388Ia2jiLw5PzNEmHiWYOyiy6Sfq8GLihe9PQj
pQ1U1+X87tRCWiAJaMAambYCwxbkQL8PQbZuGIpssxGj6fjczQ64qFwmcMoUBWBo
lF6sE8q8nMrxMYoPnRP0HSJ+uiB13ZqRHYf9pbcll+g/oCj/Nu0SB4WZKEbEy+lD
xI1KAk9EdszBQMKuTZLKR4WNeuWmnhGwLipux6KLVJiKR60B5qO0x6VZ/BYgGyYR
jR/cJlLXq2cl1seYPANCYSGFyfAAs67Q/ejJswxAtuv7v3Y3wL/Kxo76w7OpXSy5
B3F5AT30jToqjewAAbV8Asuf3w6IrtTDwzFzjf/IEaScUDSNR65YIn4s698pJVJC
X74mRqX9aweEgzsCdNJJCfEMZvZ0dc9cQY3ieLkHcMZ9uegVPUzDdw62Jqc8my45
EpNErvqrL8qfj1rJ9ewbxjx5xIvYw99y9zpiW7Add+LBVdM3ptUNre/Wp5qXEKkT
0qS1unW+Ty3o7Xw7+H3mETiE/pNeFDgErBf9K/gUvFIKeYrXqOV6e/Iw+1XMQ/tw
mEE55jNKMH5+6Fb7GPZv4/UKVyW47mCdsOixVaXNwDgiy9bBxTLN/BGE/26Wdqlh
WYfGIjxOxDpDsicgIiqvi/I9LMfVZLPtaGFimBLnrUVREP5+XRlMsYm0wecdJiah
lk422JKm/x1XoXuFMNmT3S9I7LWtbhJJl64cQFIKp3GztapdaDfAW/gIuHSc4HDs
NWjneZBQdbnXjo66DWZALn8Yi0fssL7G/2CvfCgKXw9xMMf+Bs4bVUZuxpO6KiNQ
68WrYZBBDT8v/Ck6YDQ16tNF2Tl3du/RiU0QfSsz+y6eG8SU481NE1MPBaeZ1Kgw
dR2ws66Z/kpdgY2e82UbloAbntiqOib+xmqQbaoLaSaKxhKKSHxxC+uy3crD6TFn
Yz75lIspyOT21a24Lydw59KclnxbmX2wufuhqhPbdNfiHbKhDadGoaHuku51TfMl
osXRWF1ClWCYcitDMNYaz5joGVrGCyYv2f2bM+WY6AU21DCaeCTM8LFTQoKOkTUv
purk7CKc0+MBiQxdgr+48z8KG8t0nA5AezIIL/tQJ6XFf92vs35o/DFLJmTWM/ee
xWZ0JXadtxGtFcx89E8ST3HhBx8LHFQIEyS38nXnF8Hfq/5wLIbcXhmSGEP9AtVI
rANDyv9J8MPDkyahIFNc3iGvLebub/RKURQTPsRBhjtUkV4dFDoQ0sUPOYzDPvN6
/M4bun4Q2m+BrZk/x38zI1Xxrp1GwxJTpM41P9AOfNP4ChCJKuBhqWzrC6F3SuB6
TJ6Nn0rlIn/NE6vb2LLUi9X1O6JkluCl0t3H83RgKamijkhJNnegS3ih0jTg02R6
O8kWmo6ZcXV0DyStX6NmXcKnfT0R+3SEcaLYrGNu/zsEyaaHfqlod77+sG7m9sdM
As+MBRok44Q3AtGhHRMaYvTzOJ1/xcYD55p+FebY2BJGE9tLY5FUMxu/atZdpzgi
Wsbhi72iLBA+ROdBeU3LQih8RIQoWL/E3nNnEK9fC2zZRTSu1qbz/+lJOCr1nbVK
z+XbpQxHP6Ezlp5yxvZM9mq3tVn84oUns8SoPDunwWRk3hrxnR0Dthj/Nwx7IZts
sCen15b2BDpNjJPPO5WGAsVdmpvo54NpD3b81Cxi/eh3JTQKYsuF0xV0CCtzLk+G
CMSwSaE1lF9tQLCZGWeqyqBHA+xNp0YLVMzAJCaseCdPWLWTK0S1QjK5j4qzCkia
ypFIa9FWq7nNmCQ7yWgJN+SMjTiv9caPxICSb/iSuOz2PzVVm9NMjFtqNd3YP+8D
u73rFVFjrZ4x9SSvjvLDsixxDYSq7lL/7nWchKr9NZ0xLJ7XkYGWhWXRnSM38JQC
GEyoU0tYld/qPKwqrEwgnX3Nf2T/eQXK3CfBZ+NqNCYQv1ej64UFB69NDpBPIDF+
dX50hQPXz4NxJPB7NFOou/YDHS7BC3aAXqnVBVDIj/36Qwn9kt3zbW0PEJbIvrv/
K3/+cbQgctwU0ZR1PsALwf2LLg6a9kPswRiw4Bg7ATB4c++kwVsgbwAE0VTfcgxh
xDLb4jDHEPVjSQSxVqoIXzC7TWwjJftpXsE08ubpHXcVpTmpmh/DaYVDwitRbTBA
8NsmyRGRS+AZQBY+LPxiR9FJRsjE9n3/7IFBl21Z+nV/JKR5lImdiERmEiW3L/ft
rlF0+9BTYi3DHYI7sz9KhF6i8rkHP0bV6KF6uzHZo4n2HYYbdSIt8RGSnyUuujsc
Ptv4Wgxx2ouv0NWWoxxbYzLcVyiiquxs3CtCq+wlgS939EwnQckJUyMOPiLhW6g9
d94ix00U9oOEh3+uISSVPTIlT1zh/POFfr5vOYGgvrBGNqJejw1ZAtfva8fYttD7
KLhdjACOBuKG8wQ7i37Hhe0ELyb+rFbVoRJD5v8mbs6xrdpTXDaAcf97JARqJm7O
ZXDgsDBh1O97tZ9kaq4n8RI0kRm8xid/6DUhGBmr7xz3Ac4f9Jo6hz8Nf2+PyY4o
/QOSt75S466mpAuOcWdJ6Y3ZBq9glcOEPy86Wx/p5dWV32bCInLeE03qYaYPRQR6
ZpYmgiBlIbX4pMVkEV4NzynqyEGssq7w9pV9d69jitxLUc5RbnPR6dlNZ+c0xz+V
EGATuHNE/BcQpirh4syiZczVhKzfPk0kq+oC37J1eSVL1NX13EcfhZXWRF6jpd9g
RGIxWeSm0X6ABlQ7GAEiOd/9BY+83wl+o+sxp7nOvBe+CVhpMJGkMxk8BtVIB9iz
rokP6vtq3n/GPdzXjQ19kSFF8lhVht9ihEHM0fLQZaAvYFAaG//LLvErsfOlsfhV
l75PMD5TS+7+LNxUGHmcxH0ytA528jcdnmWQC3CmSb8VQP2nhzNF/q0XFyD445YS
U/nRosx6UPygMKSdn0XyOXVlb9x0N+DFn4ymvrYMMEEEhfjLC8Q3EG3j257FT0gA
hdowCdpH+YNLWKs6IYg0w4acYDT+vIAwqUaVJpierUpgZVy+925vxM9z5lp04DXJ
XaBNDxgh7O8JDU0S0WpelWs4P77ufUUvM0JnOdam/wuFnJHydFEcZeQqoBwwXlT/
dqyPv563nZeg9AT9IVyI84MndedmFVM7I+wBjBCPPvj+KhBK73dvuUBe39OMvcGH
s6h6QAl4K/QArHmOczaDnt/RSweTFmIVstCn7b7szuZoW+DpM0InmUJ1bwud7Vgl
YLgWhzYxZk/8+tBG/5H3u+azIhMOWLr3nNTy/6kui+YFI2STt2VE+KmcJngrdIcL
DA82ROK+B7AsTwXFBefTqcL5u0l+awvxxgUGT9Q30DDL2PzK/rdLmMiOiY7SgV5w
VDJHEL5QVHtKC6dFeQjSEIzd3jVCdhhBgkz+YRuYM5oGKmAYggQBH04O8D4BFpQM
YV8am+xPFU8oUGg1xcHKk/SxB9wLdjquJOLBBAVUab8wHVtBpzcXw3vjYJgY7U+W
MHKNiblRAcxHTc811LYrgNciqQ2mTM9PGE76a39dlVX29dobNXzrU6G7GshAclNz
+8nPkSkaSUsDfoeObhUmlyN6bCwgFZXyAqKneLyRsblRZe2ArhwYjEykUAeW1PKg
h7bXtWzq1hAze122Bksxj2W569NmKJIl83nXNb7O1WQrPsMBBtDMuyZoEhpWTgTV
2f05IkECvM/DkdpBUnGJWDXgr8Rc7VLzx7UCQ+OO4yYkT4KSkdt7Z+1Q8jAS69hV
ho0MaqtGNavm9dndTbBBh7sQEu/ssDNi15Ue17zndNrIkzyDmqly0i8WirijuuWL
iephfTLo0B9zNwerAPY8lZhxCHMUii0FWjChn0nFcx0NLI45xFrZo2uJ5jjdVLPT
+Ve8N2NbtWTVFdRTXi3tY7FnBZSckVa8dPYmFPjrpUTm4Wjd5e5ctzDIVmTuuGKt
zKKKSVGLKJGT1A3vcT03HZzTA3Ox/3rcuzTK3MGWZ5OGe82CddplpGwwQXD1VRXw
CSIBIAHeiRDj7N6Ex+447eZEgnNLOqPQ9kwTxAvhO5uMquhi/R2bWXOys9oj1kTM
RVLfGFjA6xLD7jj/g3e9qqEf57dVSQlN1PnLYjv8M6NIUZOVEcJO472yjTaV8f15
TIs6b93j8sACXgsBqPk6C37Rz3cdyet8tpZtWLE8+5Q90ZjHMAenGeoCim67X8fu
CJZVvwy0MOZISK1oTYf6F0/WQBbHN0Lfrjw7hI2NfC2mvbR2VjqGjyZylHoHKHVY
DqrPKW5RgfEtgtWGzDzd/Cjo/FegCx43ED/0BK4RdpCJBDQ7I5rcgFzgIlVL2ROZ
svdUVyHy0UIxY+A/ImQXJwZMMjswRohV9/lA8gY2vuUycrOuoGpQKtGD3fihA44b
hU/T94yMLk6HiaH7209/y9oi6OL9mR/k+oLh4qoTQbDG0zPxzOvs79n3pJdnravw
`pragma protect end_protected
