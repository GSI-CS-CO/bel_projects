
module arria10_scu4_lvds_obuf (
	din,
	pad_out,
	pad_out_b);	

	input	[0:0]	din;
	output	[0:0]	pad_out;
	output	[0:0]	pad_out_b;
endmodule
