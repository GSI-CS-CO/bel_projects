
module sys_pll10 (
	locked,
	outclk_0,
	outclk_1,
	outclk_2,
	outclk_3,
	outclk_4,
	refclk,
	rst);	

	output		locked;
	output		outclk_0;
	output		outclk_1;
	output		outclk_2;
	output		outclk_3;
	output		outclk_4;
	input		refclk;
	input		rst;
endmodule
