
module dmtd_pll10 (
	rst,
	refclk,
	locked,
	outclk_0);	

	input		rst;
	input		refclk;
	output		locked;
	output		outclk_0;
endmodule
