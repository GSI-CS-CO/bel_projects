-- megafunction wizard: %Arria V Transceiver Native PHY v12.1%
-- GENERATION: XML
-- dummy_phy.vhd

-- Generated using ACDS version 12.1sp1 243 at 2013.06.14.10:35:42

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity dummy_phy is
	port (
		pll_powerdown           : in  std_logic_vector(2 downto 0)   := (others => '0'); --           pll_powerdown.pll_powerdown
		tx_analogreset          : in  std_logic_vector(2 downto 0)   := (others => '0'); --          tx_analogreset.tx_analogreset
		tx_digitalreset         : in  std_logic_vector(2 downto 0)   := (others => '0'); --         tx_digitalreset.tx_digitalreset
		tx_pll_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           tx_pll_refclk.tx_pll_refclk
		tx_serial_data          : out std_logic_vector(2 downto 0);                      --          tx_serial_data.tx_serial_data
		pll_locked              : out std_logic_vector(2 downto 0);                      --              pll_locked.pll_locked
		rx_analogreset          : in  std_logic_vector(2 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(2 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(2 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_seriallpbken         : in  std_logic_vector(2 downto 0)   := (others => '0'); --         rx_seriallpbken.rx_seriallpbken
		tx_std_coreclkin        : in  std_logic_vector(2 downto 0)   := (others => '0'); --        tx_std_coreclkin.tx_std_coreclkin
		rx_std_coreclkin        : in  std_logic_vector(2 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		tx_std_clkout           : out std_logic_vector(2 downto 0);                      --           tx_std_clkout.tx_std_clkout
		rx_std_clkout           : out std_logic_vector(2 downto 0);                      --           rx_std_clkout.rx_std_clkout
		tx_cal_busy             : out std_logic_vector(2 downto 0);                      --             tx_cal_busy.tx_cal_busy
		rx_cal_busy             : out std_logic_vector(2 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(419 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(275 downto 0);                    --      reconfig_from_xcvr.reconfig_from_xcvr
		tx_parallel_data        : in  std_logic_vector(29 downto 0)  := (others => '0'); --        tx_parallel_data.tx_parallel_data
		unused_tx_parallel_data : in  std_logic_vector(101 downto 0) := (others => '0'); -- unused_tx_parallel_data.unused_tx_parallel_data
		rx_parallel_data        : out std_logic_vector(29 downto 0);                     --        rx_parallel_data.rx_parallel_data
		unused_rx_parallel_data : out std_logic_vector(161 downto 0)                     -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity dummy_phy;

architecture rtl of dummy_phy is
	component altera_xcvr_native_av is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 0;
			data_path_select                : string  := "pma_direct";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 80;
			tx_pma_clk_div                  : integer := 1;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pma_bonding_mode                : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0
		);
		port (
			pll_powerdown             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_serial_data            : out std_logic_vector(2 downto 0);                      -- tx_serial_data
			pll_locked                : out std_logic_vector(2 downto 0);                      -- pll_locked
			rx_analogreset            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_seriallpbken           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_seriallpbken
			tx_std_coreclkin          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			rx_std_coreclkin          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(2 downto 0);                      -- tx_std_clkout
			rx_std_clkout             : out std_logic_vector(2 downto 0);                      -- rx_std_clkout
			tx_cal_busy               : out std_logic_vector(2 downto 0);                      -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(2 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(419 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(275 downto 0);                    -- reconfig_from_xcvr
			tx_parallel_data          : in  std_logic_vector(131 downto 0) := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(191 downto 0);                    -- unused_rx_parallel_data
			tx_pma_clkout             : out std_logic_vector(2 downto 0);                      -- tx_pma_clkout
			tx_pma_parallel_data      : in  std_logic_vector(239 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			ext_pll_clk               : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_pma_clkout             : out std_logic_vector(2 downto 0);                      -- rx_pma_clkout
			rx_pma_parallel_data      : out std_logic_vector(239 downto 0);                    -- rx_pma_parallel_data
			rx_clkslip                : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_clklow                 : out std_logic_vector(2 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(2 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_is_lockedtoref         : out std_logic_vector(2 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(2 downto 0);                      -- rx_is_lockedtodata
			rx_signaldetect           : out std_logic_vector(2 downto 0);                      -- rx_signaldetect
			tx_std_pcfifo_full        : out std_logic_vector(2 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(2 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(2 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(2 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(2 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(2 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(2 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(14 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(14 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(2 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_polinv             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_std_elecidle           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(2 downto 0)                       -- rx_std_signaldetect
		);
	end component altera_xcvr_native_av;

	signal dummy_phy_inst_rx_parallel_data : std_logic_vector(191 downto 0); -- port fragment

begin

	dummy_phy_inst : component altera_xcvr_native_av
		generic map (
			tx_enable                       => 1,
			rx_enable                       => 1,
			enable_std                      => 1,
			data_path_select                => "standard",
			channels                        => 3,
			bonded_mode                     => "non_bonded",
			data_rate                       => "1250 Mbps",
			pma_width                       => 10,
			tx_pma_clk_div                  => 1,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 0,
			pll_data_rate                   => "1250 Mbps",
			pll_type                        => "CMU",
			pma_bonding_mode                => "x1",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "62.5 MHz",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "62.5 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 0,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 10,
			std_low_latency_bypass_enable   => 0,
			std_tx_pcfifo_mode              => "low_latency",
			std_rx_pcfifo_mode              => "low_latency",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 10,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 0,
			std_rx_byte_deser_enable        => 0,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 0,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "bit_slip",
			std_rx_word_aligner_pattern_len => 7,
			std_rx_word_aligner_pattern     => "0000000000",
			std_rx_word_aligner_rknumber    => 3,
			std_rx_word_aligner_renumber    => 3,
			std_rx_word_aligner_rgnumber    => 3,
			std_rx_run_length_val           => 31,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 0,
			std_rx_polinv_enable            => 0
		)
		port map (
			pll_powerdown                    => pll_powerdown,                                                                                                                                                                                                                                      --      pll_powerdown.pll_powerdown
			tx_analogreset                   => tx_analogreset,                                                                                                                                                                                                                                     --     tx_analogreset.tx_analogreset
			tx_digitalreset                  => tx_digitalreset,                                                                                                                                                                                                                                    --    tx_digitalreset.tx_digitalreset
			tx_pll_refclk                    => tx_pll_refclk,                                                                                                                                                                                                                                      --      tx_pll_refclk.tx_pll_refclk
			tx_serial_data                   => tx_serial_data,                                                                                                                                                                                                                                     --     tx_serial_data.tx_serial_data
			pll_locked                       => pll_locked,                                                                                                                                                                                                                                         --         pll_locked.pll_locked
			rx_analogreset                   => rx_analogreset,                                                                                                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset                  => rx_digitalreset,                                                                                                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk                    => rx_cdr_refclk,                                                                                                                                                                                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data                   => rx_serial_data,                                                                                                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_seriallpbken                  => rx_seriallpbken,                                                                                                                                                                                                                                    --    rx_seriallpbken.rx_seriallpbken
			tx_std_coreclkin                 => tx_std_coreclkin,                                                                                                                                                                                                                                   --   tx_std_coreclkin.tx_std_coreclkin
			rx_std_coreclkin                 => rx_std_coreclkin,                                                                                                                                                                                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			tx_std_clkout                    => tx_std_clkout,                                                                                                                                                                                                                                      --      tx_std_clkout.tx_std_clkout
			rx_std_clkout                    => rx_std_clkout,                                                                                                                                                                                                                                      --      rx_std_clkout.rx_std_clkout
			tx_cal_busy                      => tx_cal_busy,                                                                                                                                                                                                                                        --        tx_cal_busy.tx_cal_busy
			rx_cal_busy                      => rx_cal_busy,                                                                                                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr                 => reconfig_to_xcvr,                                                                                                                                                                                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr               => reconfig_from_xcvr,                                                                                                                                                                                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			tx_parallel_data(0 downto 0)     => tx_parallel_data(0 downto 0),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(1 downto 1)     => tx_parallel_data(1 downto 1),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(2 downto 2)     => tx_parallel_data(2 downto 2),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(3 downto 3)     => tx_parallel_data(3 downto 3),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(4 downto 4)     => tx_parallel_data(4 downto 4),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(5 downto 5)     => tx_parallel_data(5 downto 5),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(6 downto 6)     => tx_parallel_data(6 downto 6),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(7 downto 7)     => tx_parallel_data(7 downto 7),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(8 downto 8)     => tx_parallel_data(8 downto 8),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(9 downto 9)     => tx_parallel_data(9 downto 9),                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(10 downto 10)   => unused_tx_parallel_data(0 downto 0),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(11 downto 11)   => unused_tx_parallel_data(1 downto 1),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(12 downto 12)   => unused_tx_parallel_data(2 downto 2),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(13 downto 13)   => unused_tx_parallel_data(3 downto 3),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(14 downto 14)   => unused_tx_parallel_data(4 downto 4),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(15 downto 15)   => unused_tx_parallel_data(5 downto 5),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(16 downto 16)   => unused_tx_parallel_data(6 downto 6),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(17 downto 17)   => unused_tx_parallel_data(7 downto 7),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(18 downto 18)   => unused_tx_parallel_data(8 downto 8),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(19 downto 19)   => unused_tx_parallel_data(9 downto 9),                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(20 downto 20)   => unused_tx_parallel_data(10 downto 10),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(21 downto 21)   => unused_tx_parallel_data(11 downto 11),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(22 downto 22)   => unused_tx_parallel_data(12 downto 12),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(23 downto 23)   => unused_tx_parallel_data(13 downto 13),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(24 downto 24)   => unused_tx_parallel_data(14 downto 14),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(25 downto 25)   => unused_tx_parallel_data(15 downto 15),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(26 downto 26)   => unused_tx_parallel_data(16 downto 16),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(27 downto 27)   => unused_tx_parallel_data(17 downto 17),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(28 downto 28)   => unused_tx_parallel_data(18 downto 18),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(29 downto 29)   => unused_tx_parallel_data(19 downto 19),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(30 downto 30)   => unused_tx_parallel_data(20 downto 20),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(31 downto 31)   => unused_tx_parallel_data(21 downto 21),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(32 downto 32)   => unused_tx_parallel_data(22 downto 22),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(33 downto 33)   => unused_tx_parallel_data(23 downto 23),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(34 downto 34)   => unused_tx_parallel_data(24 downto 24),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(35 downto 35)   => unused_tx_parallel_data(25 downto 25),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(36 downto 36)   => unused_tx_parallel_data(26 downto 26),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(37 downto 37)   => unused_tx_parallel_data(27 downto 27),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(38 downto 38)   => unused_tx_parallel_data(28 downto 28),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(39 downto 39)   => unused_tx_parallel_data(29 downto 29),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(40 downto 40)   => unused_tx_parallel_data(30 downto 30),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(41 downto 41)   => unused_tx_parallel_data(31 downto 31),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(42 downto 42)   => unused_tx_parallel_data(32 downto 32),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(43 downto 43)   => unused_tx_parallel_data(33 downto 33),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(44 downto 44)   => tx_parallel_data(10 downto 10),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(45 downto 45)   => tx_parallel_data(11 downto 11),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(46 downto 46)   => tx_parallel_data(12 downto 12),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(47 downto 47)   => tx_parallel_data(13 downto 13),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(48 downto 48)   => tx_parallel_data(14 downto 14),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(49 downto 49)   => tx_parallel_data(15 downto 15),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(50 downto 50)   => tx_parallel_data(16 downto 16),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(51 downto 51)   => tx_parallel_data(17 downto 17),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(52 downto 52)   => tx_parallel_data(18 downto 18),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(53 downto 53)   => tx_parallel_data(19 downto 19),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(54 downto 54)   => unused_tx_parallel_data(34 downto 34),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(55 downto 55)   => unused_tx_parallel_data(35 downto 35),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(56 downto 56)   => unused_tx_parallel_data(36 downto 36),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(57 downto 57)   => unused_tx_parallel_data(37 downto 37),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(58 downto 58)   => unused_tx_parallel_data(38 downto 38),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(59 downto 59)   => unused_tx_parallel_data(39 downto 39),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(60 downto 60)   => unused_tx_parallel_data(40 downto 40),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(61 downto 61)   => unused_tx_parallel_data(41 downto 41),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(62 downto 62)   => unused_tx_parallel_data(42 downto 42),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(63 downto 63)   => unused_tx_parallel_data(43 downto 43),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(64 downto 64)   => unused_tx_parallel_data(44 downto 44),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(65 downto 65)   => unused_tx_parallel_data(45 downto 45),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(66 downto 66)   => unused_tx_parallel_data(46 downto 46),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(67 downto 67)   => unused_tx_parallel_data(47 downto 47),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(68 downto 68)   => unused_tx_parallel_data(48 downto 48),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(69 downto 69)   => unused_tx_parallel_data(49 downto 49),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(70 downto 70)   => unused_tx_parallel_data(50 downto 50),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(71 downto 71)   => unused_tx_parallel_data(51 downto 51),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(72 downto 72)   => unused_tx_parallel_data(52 downto 52),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(73 downto 73)   => unused_tx_parallel_data(53 downto 53),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(74 downto 74)   => unused_tx_parallel_data(54 downto 54),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(75 downto 75)   => unused_tx_parallel_data(55 downto 55),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(76 downto 76)   => unused_tx_parallel_data(56 downto 56),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(77 downto 77)   => unused_tx_parallel_data(57 downto 57),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(78 downto 78)   => unused_tx_parallel_data(58 downto 58),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(79 downto 79)   => unused_tx_parallel_data(59 downto 59),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(80 downto 80)   => unused_tx_parallel_data(60 downto 60),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(81 downto 81)   => unused_tx_parallel_data(61 downto 61),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(82 downto 82)   => unused_tx_parallel_data(62 downto 62),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(83 downto 83)   => unused_tx_parallel_data(63 downto 63),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(84 downto 84)   => unused_tx_parallel_data(64 downto 64),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(85 downto 85)   => unused_tx_parallel_data(65 downto 65),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(86 downto 86)   => unused_tx_parallel_data(66 downto 66),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(87 downto 87)   => unused_tx_parallel_data(67 downto 67),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(88 downto 88)   => tx_parallel_data(20 downto 20),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(89 downto 89)   => tx_parallel_data(21 downto 21),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(90 downto 90)   => tx_parallel_data(22 downto 22),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(91 downto 91)   => tx_parallel_data(23 downto 23),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(92 downto 92)   => tx_parallel_data(24 downto 24),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(93 downto 93)   => tx_parallel_data(25 downto 25),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(94 downto 94)   => tx_parallel_data(26 downto 26),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(95 downto 95)   => tx_parallel_data(27 downto 27),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(96 downto 96)   => tx_parallel_data(28 downto 28),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(97 downto 97)   => tx_parallel_data(29 downto 29),                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(98 downto 98)   => unused_tx_parallel_data(68 downto 68),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(99 downto 99)   => unused_tx_parallel_data(69 downto 69),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(100 downto 100) => unused_tx_parallel_data(70 downto 70),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(101 downto 101) => unused_tx_parallel_data(71 downto 71),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(102 downto 102) => unused_tx_parallel_data(72 downto 72),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(103 downto 103) => unused_tx_parallel_data(73 downto 73),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(104 downto 104) => unused_tx_parallel_data(74 downto 74),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(105 downto 105) => unused_tx_parallel_data(75 downto 75),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(106 downto 106) => unused_tx_parallel_data(76 downto 76),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(107 downto 107) => unused_tx_parallel_data(77 downto 77),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(108 downto 108) => unused_tx_parallel_data(78 downto 78),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(109 downto 109) => unused_tx_parallel_data(79 downto 79),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(110 downto 110) => unused_tx_parallel_data(80 downto 80),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(111 downto 111) => unused_tx_parallel_data(81 downto 81),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(112 downto 112) => unused_tx_parallel_data(82 downto 82),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(113 downto 113) => unused_tx_parallel_data(83 downto 83),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(114 downto 114) => unused_tx_parallel_data(84 downto 84),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(115 downto 115) => unused_tx_parallel_data(85 downto 85),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(116 downto 116) => unused_tx_parallel_data(86 downto 86),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(117 downto 117) => unused_tx_parallel_data(87 downto 87),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(118 downto 118) => unused_tx_parallel_data(88 downto 88),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(119 downto 119) => unused_tx_parallel_data(89 downto 89),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(120 downto 120) => unused_tx_parallel_data(90 downto 90),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(121 downto 121) => unused_tx_parallel_data(91 downto 91),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(122 downto 122) => unused_tx_parallel_data(92 downto 92),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(123 downto 123) => unused_tx_parallel_data(93 downto 93),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(124 downto 124) => unused_tx_parallel_data(94 downto 94),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(125 downto 125) => unused_tx_parallel_data(95 downto 95),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(126 downto 126) => unused_tx_parallel_data(96 downto 96),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(127 downto 127) => unused_tx_parallel_data(97 downto 97),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(128 downto 128) => unused_tx_parallel_data(98 downto 98),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(129 downto 129) => unused_tx_parallel_data(99 downto 99),                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(130 downto 130) => unused_tx_parallel_data(100 downto 100),                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(131 downto 131) => unused_tx_parallel_data(101 downto 101),                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			rx_parallel_data                 => dummy_phy_inst_rx_parallel_data,                                                                                                                                                                                                                    --   rx_parallel_data.rx_parallel_data
			tx_pma_clkout                    => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_parallel_data             => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			ext_pll_clk                      => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_pma_clkout                    => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_parallel_data             => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_clkslip                       => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_clklow                        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_fref                          => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_set_locktodata                => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_set_locktoref                 => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_is_lockedtoref                => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_is_lockedtodata               => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_signaldetect                  => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full               => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty              => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full               => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty              => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_byteorder_ena             => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_byteorder_flag            => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_full               => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty              => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign           => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_wa_a1a2size               => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_std_bitslipboundarysel        => "000000000000000",                                                                                                                                                                                                                                  --        (terminated)
			rx_std_bitslipboundarysel        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitslip                   => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_runlength_err             => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena                => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_byterev_ena               => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_std_polinv                    => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_polinv                    => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_std_elecidle                  => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_signaldetect              => open                                                                                                                                                                                                                                                --        (terminated)
		);

	unused_rx_parallel_data <= dummy_phy_inst_rx_parallel_data(191 downto 191) & dummy_phy_inst_rx_parallel_data(190 downto 190) & dummy_phy_inst_rx_parallel_data(189 downto 189) & dummy_phy_inst_rx_parallel_data(188 downto 188) & dummy_phy_inst_rx_parallel_data(187 downto 187) & dummy_phy_inst_rx_parallel_data(186 downto 186) & dummy_phy_inst_rx_parallel_data(185 downto 185) & dummy_phy_inst_rx_parallel_data(184 downto 184) & dummy_phy_inst_rx_parallel_data(183 downto 183) & dummy_phy_inst_rx_parallel_data(182 downto 182) & dummy_phy_inst_rx_parallel_data(181 downto 181) & dummy_phy_inst_rx_parallel_data(180 downto 180) & dummy_phy_inst_rx_parallel_data(179 downto 179) & dummy_phy_inst_rx_parallel_data(178 downto 178) & dummy_phy_inst_rx_parallel_data(177 downto 177) & dummy_phy_inst_rx_parallel_data(176 downto 176) & dummy_phy_inst_rx_parallel_data(175 downto 175) & dummy_phy_inst_rx_parallel_data(174 downto 174) & dummy_phy_inst_rx_parallel_data(173 downto 173) & dummy_phy_inst_rx_parallel_data(172 downto 172) & dummy_phy_inst_rx_parallel_data(171 downto 171) & dummy_phy_inst_rx_parallel_data(170 downto 170) & dummy_phy_inst_rx_parallel_data(169 downto 169) & dummy_phy_inst_rx_parallel_data(168 downto 168) & dummy_phy_inst_rx_parallel_data(167 downto 167) & dummy_phy_inst_rx_parallel_data(166 downto 166) & dummy_phy_inst_rx_parallel_data(165 downto 165) & dummy_phy_inst_rx_parallel_data(164 downto 164) & dummy_phy_inst_rx_parallel_data(163 downto 163) & dummy_phy_inst_rx_parallel_data(162 downto 162) & dummy_phy_inst_rx_parallel_data(161 downto 161) & dummy_phy_inst_rx_parallel_data(160 downto 160) & dummy_phy_inst_rx_parallel_data(159 downto 159) & dummy_phy_inst_rx_parallel_data(158 downto 158) & dummy_phy_inst_rx_parallel_data(157 downto 157) & dummy_phy_inst_rx_parallel_data(156 downto 156) & dummy_phy_inst_rx_parallel_data(155 downto 155) & dummy_phy_inst_rx_parallel_data(154 downto 154) & dummy_phy_inst_rx_parallel_data(153 downto 153) & dummy_phy_inst_rx_parallel_data(152 downto 152) & dummy_phy_inst_rx_parallel_data(151 downto 151) & dummy_phy_inst_rx_parallel_data(150 downto 150) & dummy_phy_inst_rx_parallel_data(149 downto 149) & dummy_phy_inst_rx_parallel_data(148 downto 148) & dummy_phy_inst_rx_parallel_data(147 downto 147) & dummy_phy_inst_rx_parallel_data(146 downto 146) & dummy_phy_inst_rx_parallel_data(145 downto 145) & dummy_phy_inst_rx_parallel_data(144 downto 144) & dummy_phy_inst_rx_parallel_data(143 downto 143) & dummy_phy_inst_rx_parallel_data(142 downto 142) & dummy_phy_inst_rx_parallel_data(141 downto 141) & dummy_phy_inst_rx_parallel_data(140 downto 140) & dummy_phy_inst_rx_parallel_data(139 downto 139) & dummy_phy_inst_rx_parallel_data(138 downto 138) & dummy_phy_inst_rx_parallel_data(127 downto 127) & dummy_phy_inst_rx_parallel_data(126 downto 126) & dummy_phy_inst_rx_parallel_data(125 downto 125) & dummy_phy_inst_rx_parallel_data(124 downto 124) & dummy_phy_inst_rx_parallel_data(123 downto 123) & dummy_phy_inst_rx_parallel_data(122 downto 122) & dummy_phy_inst_rx_parallel_data(121 downto 121) & dummy_phy_inst_rx_parallel_data(120 downto 120) & dummy_phy_inst_rx_parallel_data(119 downto 119) & dummy_phy_inst_rx_parallel_data(118 downto 118) & dummy_phy_inst_rx_parallel_data(117 downto 117) & dummy_phy_inst_rx_parallel_data(116 downto 116) & dummy_phy_inst_rx_parallel_data(115 downto 115) & dummy_phy_inst_rx_parallel_data(114 downto 114) & dummy_phy_inst_rx_parallel_data(113 downto 113) & dummy_phy_inst_rx_parallel_data(112 downto 112) & dummy_phy_inst_rx_parallel_data(111 downto 111) & dummy_phy_inst_rx_parallel_data(110 downto 110) & dummy_phy_inst_rx_parallel_data(109 downto 109) & dummy_phy_inst_rx_parallel_data(108 downto 108) & dummy_phy_inst_rx_parallel_data(107 downto 107) & dummy_phy_inst_rx_parallel_data(106 downto 106) & dummy_phy_inst_rx_parallel_data(105 downto 105) & dummy_phy_inst_rx_parallel_data(104 downto 104) & dummy_phy_inst_rx_parallel_data(103 downto 103) & dummy_phy_inst_rx_parallel_data(102 downto 102) & dummy_phy_inst_rx_parallel_data(101 downto 101) & dummy_phy_inst_rx_parallel_data(100 downto 100) & dummy_phy_inst_rx_parallel_data(99 downto 99) & dummy_phy_inst_rx_parallel_data(98 downto 98) & dummy_phy_inst_rx_parallel_data(97 downto 97) & dummy_phy_inst_rx_parallel_data(96 downto 96) & dummy_phy_inst_rx_parallel_data(95 downto 95) & dummy_phy_inst_rx_parallel_data(94 downto 94) & dummy_phy_inst_rx_parallel_data(93 downto 93) & dummy_phy_inst_rx_parallel_data(92 downto 92) & dummy_phy_inst_rx_parallel_data(91 downto 91) & dummy_phy_inst_rx_parallel_data(90 downto 90) & dummy_phy_inst_rx_parallel_data(89 downto 89) & dummy_phy_inst_rx_parallel_data(88 downto 88) & dummy_phy_inst_rx_parallel_data(87 downto 87) & dummy_phy_inst_rx_parallel_data(86 downto 86) & dummy_phy_inst_rx_parallel_data(85 downto 85) & dummy_phy_inst_rx_parallel_data(84 downto 84) & dummy_phy_inst_rx_parallel_data(83 downto 83) & dummy_phy_inst_rx_parallel_data(82 downto 82) & dummy_phy_inst_rx_parallel_data(81 downto 81) & dummy_phy_inst_rx_parallel_data(80 downto 80) & dummy_phy_inst_rx_parallel_data(79 downto 79) & dummy_phy_inst_rx_parallel_data(78 downto 78) & dummy_phy_inst_rx_parallel_data(77 downto 77) & dummy_phy_inst_rx_parallel_data(76 downto 76) & dummy_phy_inst_rx_parallel_data(75 downto 75) & dummy_phy_inst_rx_parallel_data(74 downto 74) & dummy_phy_inst_rx_parallel_data(63 downto 63) & dummy_phy_inst_rx_parallel_data(62 downto 62) & dummy_phy_inst_rx_parallel_data(61 downto 61) & dummy_phy_inst_rx_parallel_data(60 downto 60) & dummy_phy_inst_rx_parallel_data(59 downto 59) & dummy_phy_inst_rx_parallel_data(58 downto 58) & dummy_phy_inst_rx_parallel_data(57 downto 57) & dummy_phy_inst_rx_parallel_data(56 downto 56) & dummy_phy_inst_rx_parallel_data(55 downto 55) & dummy_phy_inst_rx_parallel_data(54 downto 54) & dummy_phy_inst_rx_parallel_data(53 downto 53) & dummy_phy_inst_rx_parallel_data(52 downto 52) & dummy_phy_inst_rx_parallel_data(51 downto 51) & dummy_phy_inst_rx_parallel_data(50 downto 50) & dummy_phy_inst_rx_parallel_data(49 downto 49) & dummy_phy_inst_rx_parallel_data(48 downto 48) & dummy_phy_inst_rx_parallel_data(47 downto 47) & dummy_phy_inst_rx_parallel_data(46 downto 46) & dummy_phy_inst_rx_parallel_data(45 downto 45) & dummy_phy_inst_rx_parallel_data(44 downto 44) & dummy_phy_inst_rx_parallel_data(43 downto 43) & dummy_phy_inst_rx_parallel_data(42 downto 42) & dummy_phy_inst_rx_parallel_data(41 downto 41) & dummy_phy_inst_rx_parallel_data(40 downto 40) & dummy_phy_inst_rx_parallel_data(39 downto 39) & dummy_phy_inst_rx_parallel_data(38 downto 38) & dummy_phy_inst_rx_parallel_data(37 downto 37) & dummy_phy_inst_rx_parallel_data(36 downto 36) & dummy_phy_inst_rx_parallel_data(35 downto 35) & dummy_phy_inst_rx_parallel_data(34 downto 34) & dummy_phy_inst_rx_parallel_data(33 downto 33) & dummy_phy_inst_rx_parallel_data(32 downto 32) & dummy_phy_inst_rx_parallel_data(31 downto 31) & dummy_phy_inst_rx_parallel_data(30 downto 30) & dummy_phy_inst_rx_parallel_data(29 downto 29) & dummy_phy_inst_rx_parallel_data(28 downto 28) & dummy_phy_inst_rx_parallel_data(27 downto 27) & dummy_phy_inst_rx_parallel_data(26 downto 26) & dummy_phy_inst_rx_parallel_data(25 downto 25) & dummy_phy_inst_rx_parallel_data(24 downto 24) & dummy_phy_inst_rx_parallel_data(23 downto 23) & dummy_phy_inst_rx_parallel_data(22 downto 22) & dummy_phy_inst_rx_parallel_data(21 downto 21) & dummy_phy_inst_rx_parallel_data(20 downto 20) & dummy_phy_inst_rx_parallel_data(19 downto 19) & dummy_phy_inst_rx_parallel_data(18 downto 18) & dummy_phy_inst_rx_parallel_data(17 downto 17) & dummy_phy_inst_rx_parallel_data(16 downto 16) & dummy_phy_inst_rx_parallel_data(15 downto 15) & dummy_phy_inst_rx_parallel_data(14 downto 14) & dummy_phy_inst_rx_parallel_data(13 downto 13) & dummy_phy_inst_rx_parallel_data(12 downto 12) & dummy_phy_inst_rx_parallel_data(11 downto 11) & dummy_phy_inst_rx_parallel_data(10 downto 10);

	rx_parallel_data <= dummy_phy_inst_rx_parallel_data(137 downto 137) & dummy_phy_inst_rx_parallel_data(136 downto 136) & dummy_phy_inst_rx_parallel_data(135 downto 135) & dummy_phy_inst_rx_parallel_data(134 downto 134) & dummy_phy_inst_rx_parallel_data(133 downto 133) & dummy_phy_inst_rx_parallel_data(132 downto 132) & dummy_phy_inst_rx_parallel_data(131 downto 131) & dummy_phy_inst_rx_parallel_data(130 downto 130) & dummy_phy_inst_rx_parallel_data(129 downto 129) & dummy_phy_inst_rx_parallel_data(128 downto 128) & dummy_phy_inst_rx_parallel_data(73 downto 73) & dummy_phy_inst_rx_parallel_data(72 downto 72) & dummy_phy_inst_rx_parallel_data(71 downto 71) & dummy_phy_inst_rx_parallel_data(70 downto 70) & dummy_phy_inst_rx_parallel_data(69 downto 69) & dummy_phy_inst_rx_parallel_data(68 downto 68) & dummy_phy_inst_rx_parallel_data(67 downto 67) & dummy_phy_inst_rx_parallel_data(66 downto 66) & dummy_phy_inst_rx_parallel_data(65 downto 65) & dummy_phy_inst_rx_parallel_data(64 downto 64) & dummy_phy_inst_rx_parallel_data(9 downto 9) & dummy_phy_inst_rx_parallel_data(8 downto 8) & dummy_phy_inst_rx_parallel_data(7 downto 7) & dummy_phy_inst_rx_parallel_data(6 downto 6) & dummy_phy_inst_rx_parallel_data(5 downto 5) & dummy_phy_inst_rx_parallel_data(4 downto 4) & dummy_phy_inst_rx_parallel_data(3 downto 3) & dummy_phy_inst_rx_parallel_data(2 downto 2) & dummy_phy_inst_rx_parallel_data(1 downto 1) & dummy_phy_inst_rx_parallel_data(0 downto 0);

end architecture rtl; -- of dummy_phy
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2013 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_xcvr_native_av" version="12.1" >
-- Retrieval info: 	<generic name="device_family" value="Arria V" />
-- Retrieval info: 	<generic name="show_advanced_features" value="0" />
-- Retrieval info: 	<generic name="device_speedgrade" value="5_H4" />
-- Retrieval info: 	<generic name="message_level" value="error" />
-- Retrieval info: 	<generic name="tx_enable" value="1" />
-- Retrieval info: 	<generic name="rx_enable" value="1" />
-- Retrieval info: 	<generic name="enable_std" value="1" />
-- Retrieval info: 	<generic name="set_data_path_select" value="standard" />
-- Retrieval info: 	<generic name="channels" value="3" />
-- Retrieval info: 	<generic name="bonded_mode" value="non_bonded" />
-- Retrieval info: 	<generic name="enable_simple_interface" value="1" />
-- Retrieval info: 	<generic name="set_data_rate" value="1250" />
-- Retrieval info: 	<generic name="pma_direct_width" value="10" />
-- Retrieval info: 	<generic name="tx_pma_clk_div" value="1" />
-- Retrieval info: 	<generic name="pll_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="pll_external_enable" value="0" />
-- Retrieval info: 	<generic name="plls" value="1" />
-- Retrieval info: 	<generic name="pll_select" value="0" />
-- Retrieval info: 	<generic name="pll_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="cdr_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_refclk_select" value="0" />
-- Retrieval info: 	<generic name="set_cdr_refclk_freq" value="62.5 MHz" />
-- Retrieval info: 	<generic name="rx_ppm_detect_threshold" value="1000" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_clkout" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtodata" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtoref" value="0" />
-- Retrieval info: 	<generic name="enable_ports_rx_manual_cdr_mode" value="0" />
-- Retrieval info: 	<generic name="rx_clkslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_seriallpbken" value="1" />
-- Retrieval info: 	<generic name="std_protocol_hint" value="basic" />
-- Retrieval info: 	<generic name="std_pcs_pma_width" value="10" />
-- Retrieval info: 	<generic name="std_low_latency_bypass_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_pcfifo_mode" value="low_latency" />
-- Retrieval info: 	<generic name="std_rx_pcfifo_mode" value="low_latency" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_mode" value="manual" />
-- Retrieval info: 	<generic name="std_rx_byte_order_symbol_count" value="1" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pattern" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pad" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_flag" value="0" />
-- Retrieval info: 	<generic name="std_tx_byte_ser_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_deser_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_8b10b_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_8b10b_disp_ctrl_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_8b10b_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_p" value="00000" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_n" value="00000" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_mode" value="bit_slip" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern_len" value="7" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern" value="0000000000" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rknumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_renumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rgnumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_run_length_val" value="31" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_patternalign" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_a1a2size" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_runlength_err" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitrev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byterev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_polinv" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_polinv" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_elecidle" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_signaldetect" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="62.5 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_clk_network" value="x1" />
-- Retrieval info: </instance>
-- IPFS_FILES : dummy_phy.vho
-- RELATED_FILES: dummy_phy.vhd, altera_xcvr_functions.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_native_av_functions_h.sv, altera_xcvr_native_av.sv, altera_xcvr_data_adapter_av.sv
