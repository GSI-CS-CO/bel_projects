// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hO5Q3S5/5TUpkcRZGfEHaCJV3hBKwnpzlVnsM2AX5a3Ia5bY/tAtqbtedy7o3smZ
aG7naXDPaW+jErJrk7kAJHsRnIwQ4614TALZXL8ibonbg7oXlWvB9yUvx9WNMbEN
XglGAb/I0mgMGFT0Vl2M1NJgrgldJmn3qoPtzVStb/E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31728)
5Kai+fz757yXR77izD6n823Gd1utQ5iASSgUXJw/EhW3Z6yAkJUFoz5i3iT8mxpx
sO2IFOSrhgxNLPw+l4zDSxUkVvPGrypttJ5iKxJKtS5qJMYZz4bFl6JvplskaA6b
TrvmPV7eacJlLXcNOfwWpzSs1kz2WUOyZtKlb6To9eVIrdMCyEHTcswFXWXNHvns
hkCql1qZ5azdOxeoSlGe9zJvdLdTuRLKUvCleXRSpVRF8F0g/l4DC6lubJV/T/0s
GXTFIb4U2UqGCLeLL8nxxOHUrs5FzhGdxlJ4WmdHe4zPlCp5GNccFI1Hfdr30OSI
1txSZifkR4VvuE/6q6nkd0gvvCCT24o/AqbSh1DFEY+mTYI+FhH9wDb0e9VQy6Na
LJaBhsI8pmPCX4Bs+CkCMm+YaPrH/tnp+AIWdQGupWSlNfyf6o+PxPlVJZjQKob3
v8d+gxdPvqNwwQFgDSbEgRpUoIaRy70+yNIbc3Ycir0O33NsELeWFFoyr8SrEa/X
BfZPGodR+xiiIIiazblH0/VmhQ7rY8oKL+LVxeDnG50BUvazF1BtzgmYySGd7E/R
BCtojgTUCnjW2OgtzMy14zJEw5x17RHJ/HZ6pS0KK2EaOX6yXNVBVsLXYY8iC9F1
9K2BtViP59ormCYW2wru0jGc4mM7VM26ElMKL+omsiZbNCYcA1wwx4JlZUZclHvw
vUdQ6d+CTOK5P1+M/zVsQKmFDRfD05LPvxdJJIfPIpCsCEBqxaGuwg8Xhp047JEy
KaK1OXykMfKas9z19wfzHGhJNkw08NpyMJBzNnm1i2yD2FucHopFeno1QDl/H3xr
dHGUBKd/EPDSprD+MjzpwTJwJ/Siof8VyyzWl3OQIKDUtro/PY7WtQ7QQtPcvy0z
80MQlkF4S/nunnzEvTjLOQTcd+Ab3Ehfe84PpnVaeczBWSqsLLa+YgEkdNF8z9lm
rjBD1hcG0KhN/D4D2KLrV5xVyVxDzZJ1G19OIgnq50LAarmXM2ZC1BGYJKmMtATD
bKKtW0ELD/Qggp+E6K2NRbud8Pw/XNmFrN3ub5S75Qsbx/korzK9XiMjFocfkuiQ
2VkPJZjDczK3KnTQ6FKXV2kUY+emllNzteJF7su1btcuYpLlaBCFTP3DQP+zn3ZP
kow+P7ArbVTd87TNfVzMy2WYyUUk1jNfOFJ518AFXwm17t7T94704hQqKZY8k2h9
9mHgpvV+NHuDx5HN4caxPtZL2bsPM8jVlUK4y89o7e/rZslJeaBcSya+qibrzz15
7ytNMjJyh2I7wpfud252zFcxhQvFyFHZ4Ttjnj0+k6acAUvZGOOvabjmb9qtqwAn
SJ0mh/4Xvr5yZs17wY5P8xyJd0Ca1P+S2EVDMU4uwCCWmOZcdzBSVWb83zgfNhDW
FJL6WGZ7Il5AqPTuSHhcubuEDmtXudRFD0bjh6EXvVqyHfk2oUlkpNL2JiKVCHJr
6P5sbuJSD7MQHUITX7qg3in0A6hWkkl1MRZPIfGZkwOIHX+3tdbS6nl/yx5qUVbF
Tk03Fs+ZmRjv+AHqPFYYa+n9mfSxmOl+AAP68bWvqHUT5pOeV0qKXQtlSnkJCW1c
mHSo28kx4LZHNHaY3Gqkni2FjFPd/eReTLlRFWz7nwoEfiXcP3ScOP67lFvfkNtf
PL513ZiChlk7bZVI0YS/ksdZxpoz5jpMTNE+/SX4V465Hi1knZ32EUoYH1hqmM+z
0Ep0nm3JIADDtYFbdPxSIZb1UOt0lKh2jDcNsx6sHmUgUw47FWxu56A+sM3lPCuh
WVMuWblOJu/NtyyhivZgZ3AVPP/fQL1nj9wtt4kP3mlz21jkM+a12Sh9BLVZHgm8
sxH26HzdX2olCMugG2s7QjNRo5XGKeYWudZflYd5IkX9drmEUiXyeX3ap9XUT3z2
Ep5v3IvTFAdVdYgUjLTwH0VHbv//Khdkwu8NIUBswPYNpM07+aTlREqHoBBpJ+30
472XHhS3PoxrYyvqZCk51zFrtG0fw0VdL0psoPnbDf+x194q4f5rEOihwFvhLYWf
tu9fq1EVz0RjzjPvS0hvIA6Ipo9z6MGfNdlLg8gfq61Qn/XqJEMZ8y9SvcQos1XF
e3yrr0bSr/tbHJsSSMiygCVEirXBL8PlCpNi0SvDSpkd36ToblZJHbRmD71GwGhJ
6UU3wplFEbCprld5+oGXo+OWQrxSFbixJX/eBdpVHpB62+Wdy0v7hOjPcfvfPIRp
Ur4iTp+8mMp//OuSC8vI14+vVOAhX+OVkpefZLwwtnzPa4v5xJfKY2zLYZyA/9Np
tDJBU6fNrhNTAnAMpRNMsMVI52I2WeSSP7qW6WyFkg4TIy0eenYsNtHWxEfcaPHp
xW+OC3/R+PSe62Q/vB/GJ69A64n4CRqxtwXVchWi4oxbp/QPavQy7QFIlYOH8MLW
cG+jmaJj72Zse1TduxdQ6UJyKEdn13cevL6W9kmqrJ32RgunL7kxT1j6kqlbfEZX
uf8iquxfNSiuVaagv/BH3BEjdLHG5vhbzG7Ep5xkJvOce6t2m5Hnj+EsVPZFDWSv
3n0iINxa8IAaePJrhH61z07K+L15nGskFglfJ1e6HhC/oicG96GDJqj1PIr6kL8u
R/NidRPeD3m2zHdthpCOfZussxzugF8/a1BRDrioEJybVNb57OFg4ZARZNY6hiM2
5TXT11MRy/XoVFq5IARQ1Nvdq17C90uejvVRAUnhkHByEEJN9Q06IA28SWOV6Hy8
DoPfJi84dcPo/Vknrdpm3oh2UlEUbGhM+DrehEDY55j8CB1me+d3JKBhMKYSwX1Z
7I9fSIZYCyIkpJ/cIUNliWtmqUmEH+gH7z8UVTm1DTtHLZ8VUe78kBemyfsvqxl0
O2AVgqK6fAoP+ESBkmKo1v4DWQNUtEdaux+5voOs+JS3Ddwlm4yU6Vfj+8mfQjHL
N8NaivOY3OBjxwtTJxRqXz38Mb5PqFJzU4iU2tl0sCXw8Zw49auYLoCHgq6DuGrQ
iTXj7Wh/jJht4vzRMcnjn1bFtCYV3wXrX7wtzpHclOUDAi2YbtQnOLzWPwvbO7M4
wu+D8bVfxGMAFwhgTsnNNMgyZ7qteD1/peQAan9ruZlEetfbEPLQkReLoUPjNYsk
thOyCeuDuptcwBMemOoPQ7j58feO0mWc5nlLaLUm01/DHJQkBFhKnnhxIp16gti9
UGIMwCbNvR+UbYWdF8efbrm5WFIA6Y3m0ZWNzbT8qnjaxDxKH266u1JeGSFdHvEg
yRag1KdZ79O+ywP1y5hTVVLa2msyLc4S2N92JPgppWgTYFnQFq9k5vgtpJaItFsl
ynb7EVX2Xux3ZlLlZZooEqRlYRV7U3lPo3Ghb/b+GpHhO+4e4C3Dw/2T6COgaRxo
YY9XN0BQqYnG27kSvOWpebCyfGdkeldCDwnM/NiUJ9F+1rnRp1nGYtETojIQkD1l
6N2Pex+wzUfxFwAvEtvc868lxhip85X7S2eJ+AEkoSYQ6Nm2Vu4AaflzOTK4LKkY
9wIbWJY6WCetfm85Wt6j0oVbE3LqE7tba+6QT8zPEAbvbIyyl3bBb9019MQIMO8F
GgI4OjMReiSpXcEf3oVowJ3DDaFHUTm90qwev8Sg8nCHJo+ujBp5foqTJGUdiSO/
SlUrxSVVYHIZjpOrMQn9VCRhZcFJhsI1JV+HZ2Nb/6QqFr/PxTvgXnYTLyGYeVA6
dkGwvH6+tbnW5HFgm14Dl3rQDDqyDndoQtr1+UUJHCgUzrcCqHlq7tR4CxV72OiO
NhLN3q4l3ZAzO32ex5DUFfj4FGL/0fFARNzHepvk/PawwbxTdB0QWCo2KR8LIEFt
5AgpHgs7tiK1KyqrFtM/GAR3Ow4kJFMU0e8TjG8rCaqnOJ9aJXrAMxw08XCod9zg
1BmIRyNHFgkofuVuWgMHnqfBCBYbiCjvdu2zgpBNebzaSxQIJityuTY09aEcoXSf
R8u7qNIcocPKN88YpzNMcG8DdGdB93/qbRPvdJiIg3R4r9meNWZI5qk8j6UPi/Ov
atL98e3OKAvB6rItbLMYhRwIYd/aQCYSXZynR3HzevVkfke2dzBhy59TGvjMRhUj
9h+LMUXPm7n8vDcd55Jqcn/OJ15stBtSBFzscfafMb7vNy0E3Txq+s5J7msSW6Kr
VmPew2jNVZdhMkWBj4PG7YlBX4kpnbG8T+O+rda9Xpv9R+7d5+fpVrbicCJlHI72
vUN8FpZV0vUIusOC3Q2UNDAVUL9E+GXJl6nDJX7ivdAbCPd7whUcL1vObe14uMio
dstwmKeGpNj5jHhjIvl8cajO9dgrg1/AL2+5ymWZ7yjDqfm2IOkxwFTuzyTlluqL
pmgVXUX9GT9wNSqjG9JfkA2lyG5hFqaRlrtpzGX8pgTByZ8bBi3iReJvqrtUEtxC
m6U7RU54EOCtyXvEuAE6EubX3LBRI+EJUxtAERBy+QXwQqgmRXdWX8koEk9Ap9NS
ijEPYfGt9WYEZYtiEIYWNGDEyGw4WhgbA9gZWR3Y51MjjLwO0oKj8GE3kc+KvufC
PFz2+FMYSCY/5fFLv+zEbGn31Pi46JgJcZiSh95Mez227GsexBULE7DAnAa8xqtn
5aqKRQ1lPf0M9k7doIV7RDhYCNJFUkRhxkz/g9jxoMH2FVh7A2X6cNoGaFwZXKD3
DuTKEfpA85JfWro1uZwUm30aHaokPvyP8kzWE3WUnerd0ajBJVTzNCNs2l8nAhH4
Mnmc9jIUjA8zA0q+uTe4ggXhl+2jeMeNNHATMpRY5uAz50sg8SLB8lAtTmOd2sFL
eAjni+lqPB50Uv2eyOhWgKSKAv2IgdC++xhscolk3//iFkzPi+N4Kdw0Q6pNHWfy
aQLPqqt/vSy9tBZZSdc4OmvAf0v45eVB4T7l3cp2XOntTJR84lRHlASKXZv977Zd
iwrQSktRLJzRgn9k2YnyylijOP77J2kczBReOSNw2nyxQI9JqB5BWUoLkp6ZFL/O
3Yjikdishb7GlpdfOoWIx9qT7UjidLfWPwl0xfkAnlNe4TApg7xIGSWm9CCnp7S6
LdpOhJA2CPOMkX3IX+RSHPtQdlfUEkoArUlpojcCftWt+MytmlyjlhjPDQ16DabG
gGRaT/LuzTnB6pBnvfiDvO31P1jeeUmTIC1lJvrVnTP9UFG6LnV8VwQJ6pzfEdEW
Tt0VhUPe8t+Td8LmjX92uY+r3WyBxMC3UR2UWpUOLOuz0ku2LixMok3jG9Hqkje1
OwfyYtJwhvUq+OtMedhYgaGzaZcuBEiYMl9j/m4NOxvKHsezDUL2PHz9RIh0RWDo
f4c+gNPJK+N4zl6eeVZtK8R8oiPugjBYpcFt2MByVvvA+domfO6Pkf36fG23pt4c
dO6yZBcdwqTUT/2eH0VsdhVsSuUTo1/8m8evO9Gr56HQZJTCexyOefa0XnORyQg4
ZvOF0ip2d40dVTbb7sdrCZsmCJ71Dmoy8TfWiHaSCQuLHoS+XKi/JqN9Al82refS
qvDUjV58OaNgZLecIxyNT0uFhqXLmEkDZinmZNKKYctIc1K/XK+Yi18r0/KYYIM4
jcx1Pix8XtI2EbkJubHClas9kySO2GtrAwUnxqfjsEgV0RHiadyj3azJGxAKpEQW
NSBFuUw1zQOUcoWRMOkZX+P/ouctLCuOgIefiPbzspZChIkznWI+MdKS7F2EBxNY
Bt/zsvq/evgDfcX6T5r50FBzn3fx4FexTfg/Q/I2oNNrD2d5kXQvqkAWoNGC51gl
0o2CIADUg4/KNLahJqMDsib97SvfXHJmWce+cwBK53zYwqAbe4HTKgLNTzX3Yc+/
VoCnO78Vas59ZbqCUv6kZNfBo/ukqNNAzN8tbpjOCw20yUBQv66ghIBWrN1zG72/
Jh3SeX8m2HTy96JrsA14eT0lxNHkYu3+xZjH5QfMphIyFLdgd97tF5taKOtwcwVA
rk/AwHCyzakaw3srkT5HP0MPdG01vQYeVIujvro/zWHIKdvvE29EB2AwNJw8r909
2Eg38Hklm9smD45g+DSV+5cUONHS1HIP29wn2Ztn4walWv5YOYwbn7bRun9Z8DdF
NrLyMqedtXr9QYLsuiZv2NxoUQl3gDBfJz6tm1Kk57ijoSpeJ3VpaG8dxC8C4eSr
NO6+/3bjZTwuQlfuyDzUVTbm6Q1nzjQKW3fLPBCZv4oYf+zuZzAO4WAImLh8MaiJ
IcSVzTCL+x94kwXW7Ttt2czxoOIegz/7VxQQXD33bHKqFqI+C3lhVUUNK/n3DRUc
uMWOWXv6faMx5J0OMMRM4LGIhNz+2a41StdL+ufsxFEB0E4k10dpp6zG0NY1whXN
m3QSCR4ceiEWjeJ4DTVNpGIG28tUVG8hWd/pStu9NnAWeQxJ7nqwdy6AP69mKVK2
07gwS4HrbdFbrR/18i8/ei9EJs/Cy4N04dOxVCmncbUKDXNEBmgJWraIqN0aAFfD
CQG5LSfqbcWmKQGgfv9kHxBwT9ft3tQAq5ro5QltPRX00T/GOUgI+jFfXr8nhRg5
wTR3GiDxdNXYjvyxKcs0lDEiMAl8KTefshMiRlx8XnTc8LYIy5/eLbc9z/LoMsv0
XbUSnj+wV6Sm0p2G5qnwh9VdIyBC3vFo0t7hlkxcl7/rYbjVBrt4BXCOLcPYD2pS
OegNwgmBC/fzcDL6l2Xk4d5JDaDESVZuljUaOaaHvobn3s1uInQdbhRIllIWiO8c
lIg/gOT/m3W9qh6U4637RM7KRM5hX06RkgO/ByPKRCut3fxslBBuFWNCbXrQIkI3
xI6QKBNG1tphEoZMlmkcIuYEKTWiHPOQCRLo/WoMFmpUb2D6ZqJMaf7FR1vW++zk
mBkfkETR++vTtsV8FOxqlCRAt4EViNV0zegFrjlQDhK9HNJ3UEPXa85JZi7ORsSX
I/uywh7dTG4bE5DYOyYUuAVhCL0byzlCrp43KrQeTCpELtY7N2JqJolkpLAvm1Cl
cm8iCbgP9tcMDXc45ZL4Wy0xqqUTOssqIj77ki8wyNiBVKA1r5Ppdp46J/lpiytp
M50wTJjOeK9DN8DE7ohDoZ0S73rVo4+o30i/iBg+uo2J/7bISBvwY77JZKaWSYa3
dDPa6D9csAD3hTQyHY+v2Xp9O6H3R+4KwK2BE9po2Ses9giSWUexM6auxSKSzuV4
v2fpUbhkORLl19qd3MFxuYKd/UX8Uw/JPJNE8s026B5PWk0jcBcJeDceINteOXRW
MvdrsEe+j82dJbVkkeIWJxJ3Nq1WWLcEkIUlyVQ0Remwi88RnvCmwaODx/s2glsZ
ka2OZy/TgU/n1A50QCVg4eGibfjTpLOACP6SXDnv7vpqwHzqNQG3FhQiEgt7xG+R
Omw+PDAQOxFYxWGWmV5CZ/C3Ugh9t+q3t0t9quwMCgpR4U1e3/mu4NL+fkAP8hNa
HRvBQKW3annhoLtI2cINNWIp9Ctz2JErTticEpqtPGneRXP5C/yJpKanxXSsVOk+
OuRd9mV6LxTYo7Qm7rvMuoybqR+yTHnAcuO5cBDX+jxCwnVQuuOiD3xBrzjJ+tx9
CIttYLxyD45V5cJoiRsLR5B11oJmeCSoUjAqgcddkHZ26ruP0vMauLA6fQ8mFZqf
CzMgZUcGD8v8W7uS48UOy+EZy2YlG8S1bWEhQCJefaqVN5ka3MwOTp+sT+kHkUBC
jOTUA+0cn43/S6vx1UaxY9scndVYB4bY0fEps4s5uW+pibwJk2QeZDdUNl4LIp5v
Gp8hWn/qWPIc6RtLDIhLEbPUv/1A91Ty+Cf+4fyllYblof0DM7UMou8oAahKJoMh
HtriGHQi0Gwn0KY+4XJuL2mdjgVqmjM2R13V0e91aG6b3iff313Y5v5iJphFVN4h
DyhdxSx9kWOVZpJR0WQRAY6iN7N28dLMEzNALUuTviR7jsbgByQa54GQ4ymfdBQo
OifEO9MLHceR25v6RwQAhC3tEEgZ4jiLGUNzaAMfL+xkDGE1pEaA2f1VbQwmWfsD
Pg2WlCySCKVkAo9AsFmYdu0bFR9RsLqti8dIzOIQ1kpnc8gP7I2QHCMcbMa4iI2N
0FOExZxU4tuptUw/NOSAM3Vq0KB+IgYIN9LrVHqH7ig7vYHMtjPyAPVPELQjC9S5
H7iQgNx/aCov0CHgDl8VRIyRu4azq6PjQDFp/Bj6iF54vDrJvWe/KKEmN2E9yLET
siKlBCjzIuaMKABh8mwYrDteiQReYiLPtjbFEDPVMUOG5Tv+FQ1x1yMIgLpWsgP+
Bh3OTCEjE5oDY53aV6W+JAuFOfxBqRAjpGMfsAq69s009oenBFv33TS4+gizm371
sV001eCKu+0ut/9aZUILpGnK2Z8eEgrug/onJQb+w8+2JQMwQWFP5GJPKTz3jVhH
EzOBMuyAP7okjGvTJSFpR+3Wj+ByfF1DMTU6Ac7n8pIRccAxFpfWgEORuCDffjYl
06+L7UZWOR3/iqC4uMG/+tf+3orkZq+kUlhOJHsB8EMPfOcl9KDMTPTncwUtIB/U
zMENZcxQtUG5W1LObRo7xKoFcUZ9ayr2iAl0qKVmSUpK2Np+icl21Mca9IgPLP1+
XFlK8da18wMJsqxIIc6a9vGf/JSFixJkQ62Nq4Zah/G6BhxiMgJjBDDDyz9m3GFG
6JQ0YH+4JUx5WNoVNhrZAmTzcKal7Kq/22b4UVOVB7LcBPywHeoyppv4aUKdcowB
IqyrFJUM7OUXrXgDrVF4m5KKqxny94AE2iKcVScrLqiyFargmd0MyYKZ5+npE25C
SCPqCy7LcXpfuLMSDQzeFCfcg+kdXsxUHmoJgVtn8mkg93CvuWIRODHnK1Mu9/0l
JOUuOi9lHR399piuijSHalCLQ7k/tgdlhmBICZN23hReBWEesi9UBRLuDNJ5usT9
dkuPkzIOpUDvlIj4uvQVULc7z8ORIc5dojsijht4ETi/9ZapxjT/ElUVqq+ZLDFc
eOsRvnpo7a0Xc9/v906EoL7klbkYLnLzyxyv8y/DXLBcpzkUD6Lbm6UZQuj+oDDQ
H4UMj7gl0WD3+J+JoVkmp1254OD8vdOXM3GGyIpxjGMeFklHRxyd2K+1juoQ7B56
u7UnApttQvU73XVf4SLK+Txn63kACeae7QqcuazU0IEHHVRSJGoIt2y+OL696ocR
1vaH8BulRCk1PfkY646setdSXNCzRkAwJJsBNSEnRNy70s7A6acX8y+WcAzNp4Xh
TK2nP7z3A6AGWDc4e9Bo6X9cQ3TQSDT1/9XfyyrqXF0JotNnqi+MOQltXtVEjUA9
jmiuCPuwhV6YZA7pbjgyiiRI5bjfb+vP+VXB4tBDiWxAl8FEf8wFfv66Agsf3WaQ
ZCmREeZeqzT8IQkRuHQMWHx6MQ8jGQtE1KwYE3L7aDXpu8xw4G8f7f+0Zm74PMM+
rLKNaE6z7OHypD9aDdNn1db3oygdxfhuCMJn713r7tb1G4IY9kT0vLwd+BL4Po60
wMfEj5SJm8C4acQ3ZJObqqeu9LfsMVp2x351IvO9fefG/7a7acQnTidFJs48pHwR
uDT4qDTVF/312FEEIKZlbDd1rL0xRiHhgKZe3BXEyMdDoKZjb9qL33HwpMTPxL0o
20b9HXF9f9m99a8KSZwrACiY4HW/gjHdRkv5MsUxeN5M45MTkudEbuMIaxHrxv8/
P4vXyILmQ1xb/s9qZqNpC/cK3FNeWd01rTT2lbxvlNSpiFagiuwxtEGYPKCnolsN
dz2nP4oHJnyasbXlJSrqK2zIeOp5Kb6BjUghDIxKhJ72ttuvnMB032bbtfjfmJ+h
IV+HF9xvkssClzUOiYbxkY8pWQ1zGCu8UdMTZPt3ToNlMcbAVT/j4GIVA5SbLbK6
MQRHioRiGDw5HJDujfWNBg9SqQBVrHTbU831FS6bimD4vB5+ZfFa+jur/IErrd3a
mDY+xpadqYBC5/NmLa9+JlEM+y+4vyRj7u42VV/eINyes5QHCPcaWunsDxf7fn6K
Uc/KAWwNiEjI9rO0K/PbwrKo8AI+EvJdggtimtnPDpAJc8KL+84cKsj5FybTMVhn
JYZ09sC37oM0O7JbiLT7WN+tVXC9VDswsoo2Qv9HpraniyXw79lc+P7A9KH/SxAD
YuVbIHq87uhGOxRXL9E7Zmf31KBCbxBVosGJ0WZQtrvbDsgQhRcYLJzaqxRpVXiv
fI7hdTB+1hun1R2wrkYJmaBOd6yaGkdc5VhdNrs7MGSvCe8UEfHgGVN772fZdHpm
JlSKZm5Cgvvv/ctlAAWmmftXyPtQM1keJzoW9B/bqK+OOm/Y5bmeiCBKOfHVDGM7
6ZKmeKdEHBWDuEcyRMvU2Ih7RVAMrVeS6lUHvAdFbox145mL7imy5fcDMjxtD0Jv
cZN4IogbpwT5xv45hhstA6ASiIE4ajLf3sSyrCYlLITLPdOoZIPGlEA6Gw/DCnJC
ohqSoNSTwUpF93NrNku2sXAUMQ2qPaLrrcgWpFXzUmDpsV++iktdTnIHwqGREbdy
pGin6PE6P4iBd889r6GVL1Aud41Eliz1zpot9a9Hy5FrShrx240/PysrfOwqQJ58
cWQw2oasxbC4BNucwhnQCUkXTv9glycUeQVsXNaeIG+bph/d9Fr8DNEywkmIgkHc
COT7lLHwfElh0O7mk3iZlOhu42DEkDhmwXQABt1OHH4ltKPbs/LBPECrdbJ0CZbi
QTTrlze8tG3J/hHNnqjA6KcBEdZ7TXh6dab2LgGMyodg+k2GTH9n80Utt4ShFNj4
ohlyvAFcc2VS1wwArY7zR1iokn5f32IEhRpKBISHjkJgVCq4/6ivp5/cUQRG1vP2
dTAuN2dj4kA8kqzhmvgekGR2tP5HIbQbMUHRt2jXgHtTDnPNmTpRMo07MNeeWv32
e8Tjc6XoxyRAO/PqrTGWBp2orlGrIDWO0h8jsZPonue2WLYeSsEvEHqg5DJ4v+kc
/vJRdUERXBWhrJFE7tSvx2SVlcBmyTGmQ4KB8uKG7UEYXEXgQD5mPw5fgUDayARL
b6xf/ySbX7FZ7aZgsXwGv1Y5EMf+BQufJANhv8Hdg+H6xaPOL/wHbLhZiWF1vz1B
K6GdguZH3ogQWmpg4rXOd9T0mgNK7+vhhm4NZuqhsA88Z3TjUsWF3JDv3DNLUB4N
j/0y+k9URtFZK/Rfzf1a8UDA27k4ZpX+ErxFs0fSfxNoyqRwwJMTK0mZCyevK66W
0pVrJ7n0cAnrBP7bErTb1zr2LF6erN39GRdvzfekD1FgNO6ra+xBXYRRZqb/I122
HPOQ02ane9XVo91AM9ZWdvtxyn8cIfhO+p9UDjJJFcx8uMxiL0zd45KL1U3OX6r8
IUzaCx6mvf7wMJQdBIXBRLM0H30qheYNGmqw6yk6Pkp35HOhDE3tT9LyYOKfWgaN
sr5NDZkNmm0lb0AfaTR1gxj0OscPopZGYsqcsgf+oGItVSx9NsMlMqc7X2dxAW8b
ED/QstDQLFjv0xBfirLXEWSghVIa6h2j2W2h+DaJ4Nsg3sEk+nyoT/k7T3H47xBk
Fs5mjmtjOvPY7iV9hOoEDUYILi0sZShmS2rzt/gJ1+BE7cWK7eHLDbBUXP/cUyK7
vjQt1DfnglY/d6iZxzujZvI8cJndp9fX6s6Ohieh6vZj7TU497E+FE0O2wP1xXHW
v1s6doJxdkbc8Ftkle9CE/ZJNNLE0KbOgM07xibyB0/MoaBfbWfSsgjTcGxc5smd
UGd7YksLy5t1Gitksm6FjUQZBhyD7aIeFCV9v50mb5zrLuMlaP15fyhlrKBLuFNX
u81KXTXfSJgDjsjHeiM+vRGVcVz8A9nDVrKMXS7CAbM3wmeqLfywLwDmRl2FjRmB
yqlHn8MxKf7s+PbDSC6GklZHsSC1knHrLO6ZK9Kw4kd4+sPjqVS9sLPTh2zuoWMe
xWSjEBq5T9UU+WTWkuJHv/4eqaWFNM4TgF/YvRn2rbLv/ks6DnQhobb4Adj3id1M
+4pbRrYC3WYP6NMweUBBdhcUsZkkcAtEjzOAN3GLieHXcqlT9uh7AVne7KMhHc25
bGs5yqvRqUmQRG2tqiK3UcXMuTrx//LhllTWgKMHQ+MTPtxph0Hh0GNydE0hLIMX
p2M9mE8hredSg9vMPVUhtrFmLi34qqzETWRG3MkHEEVSaXJVwt4NqPZcPk7M6r/W
s7c8edVzIOJgmKakkdVwkiVgVTFhGuYI3k+b1HOIX1eXhBbka393lbHTm445PNeV
c7Ay+RoNE9PHmcGCOY9YN9LhcWQeudiNKNY7ntn1icIwVFUQ4qSDe5LndGk15nGj
U1uXZAoXdpVrbnmKaqReBSQ59Hm7xh9p4jMtXw9CCwurniaYAYlgpAM7RnpLrjjb
OBLkO2qAR9VC263igydFAqyjrGVoIcmT1sZ5Ix9H99OlwbuSZz/1XnDwjiGQIGYR
mpboX2W67axzWDA8raMpdjE5f5U9/F/n4zB/L2FVArV+ASSVZYZS/79q/HEsLd2q
+PdxNExnpUclI5tNfZMdLzzH/rZqqoh/gYCc4/pJZY/24xFQfpkhH3O4UJmq5gO/
2guVmD1PzpkC2xVtCGwzc50OWpE56BCF95YkXK1zAkSJM18hB6HBSFtXvZRZa64j
EpJ1hjkxc6nX9G94jQ/IkwU/+3RiR4wO6hHGPxW5eObIMEV2vSz8OYiuDJewU3JR
ohbQgEu9tyvM754jZmWydMoSR1uRwhxgRmWNB7NLRf4vM1MhJ9VDkV7LcazNB3dY
Id5sMQ9bzEwSCk0txUG/XB0DeNfd/URH4Kdgo9oQVTTkxaDnDRdPo05299pKIO+y
FFPKPmLMBDhppFAUAEHV9eRvA5JowScBDvl2lGML3BdyeR2kUMtyFzqOV6ey0xA/
UP5yaWoSxW2Wheh67FD453YEHSNqVfUR+vox31xlPCxAN2A+afOpZUEGT/HfWMY4
IMbFtww0W4lF++gb9QIvBhF1PuGFQDS9eQs/EZqWgOgoSWXH/x9mvXaXJ7NaYsbU
yCGHUz0DGqRejrHw01MHuqVsQGMnfeol3bwAEbEs/wbL7kBKynt84I9BhFBOuWZS
fLx39LjWpWh7fMEr1uXOCbqDKsfG3CgbyZEnToo93LRQPP965Y5YjcLH0rNI3Qf9
kYv2GV5KgLD/sTdL2ylRVpE0E0eKQqS5E+lkmj+bCu3Oa+sTLtyBpU8Q66igiRF8
TD1mh0LM9L+2o1u0byW7rLcyBQC61bvtE4m6m4xHW3MFnltZhcCWvZ6dHI6ZgKAi
Qwsi6kNR3Hm0ywX8DaZstPhaU4e0t17iZDth2JTX9U4L0vuYLLSkE2zv7GFbSeVN
kMuL2p1flZUELSxPO8p/i4DuLhYYuhRwN03BaBuiM85skLxmoGf1glJdsdmQC+QP
K1r3k1TLOjzuJME+XXOVKENaeOWKsCnlKf8ZAo+qJzr5qE+oIJwVYi/psMlBvsMK
pfciinuweYle4Yd7vQrKQqY/UtStLrczrZcoG7VQkxEmIdQRTA6rO0kyIh5K7wHM
w8icvlsJRVK+vGcXZO49KUCmw4p+ZYUleXX+sSHRZbjy9zT2SFi3eKu2E3l+RcEs
1wtI900cfUl4pEJ5fVzhZMCq6DcoPjasiGUSeADsv0X0+dTlvjhDRWoWbu3/r9+v
V2wGX6w7imIRy6U6rWmdbEbK4Q0Tl8PkZ1P3ssRzTA1Ptsonhlf18/ulNIH5hDGb
Mnb7Dd5K2Ra3f+YvVBMWA7/vJ6worqd44TcsrL6swqeN0bYRaHQ0t9drrsNh+RH/
duIfh2alap/uV4fljP/aaTbDMbJjs3d0QhUekFNLFgSQceXPjGmB9vl/Tx+Mz3Jg
iVnd1paGiMPfYiM8M7yoUUbFJR/ATUJ5MdsyVB7UspjKNt7alOzhPtxLVfThh5OX
41NvmBcYiNwOCMPQ6BswxdHRgVQnaXBfi/nqKaJPz5Z+RLhjeFs5NQhEdReWrCGA
CvqP9SxQKU3x3enPzopEYSrLsOBlIKPd6q37eg1oegNpzxwZU8vF2Kv6RC85OOYx
R804EBfb8sp7zBJIBaRa66735RlSqNYj32e8mdUamZAg9Tdjhh4Z5hqyqfJHn0T/
+wZRfhNxtym0SkYMK3IgeIfoNtYPvqAsiYaHaC8yuaD1FbuuJG0c7hWwXNwBdKr3
k8OSAsXe8SdUO8nfif5VONynckFnOhSgYsNDuNmXQeWxaOKWJNTsiEEPGeR64Yvm
YBLMCX9QS/+B6uHKa4iwD97F2MEMUjJ7rqm1slzPK6fzILq+2kgirGfO9mugxkao
vwYj8CIbXfPk2npKah6mBa4uFsnxEpO1PtlfWIQ17y08W3KvPYfbT/yMGYbQZvRz
McSGvLN6A1CxXfOJGJi4EkzdKhTjAnOO6n3EZUeOIjKGHKSoQczpQhVcHPTuOtSE
yOJFSKCMCCS4FFEAEkDUdP4g2YTvDI5xK75hgv9dgtG7+XEam+xBmjRiFF8+V0AJ
IRriWIcmhMIIa2zjU0j0Ttps6nB9I03mLroznE7N/7G7kYs9JhKPWnoYWPMrytJj
rXUvw1Hi0nRwbdrzgEnrGWsGDTQrBf4yrqe/AwVjqhVQ3cZsrrEo2gNZQrgLZbbS
eBXIAdR1O0psOqtXCCt1HshUxYLFe8tWmMeBtdupsF1tpMPdkYAHX6P/Ho31t9yV
8YqB4HVOqyEk1aQ3nUkCybPNIqIlEbsE4mxnfYOLDwbdMNxZ6VTTzQhc8wCaYy8S
d7suUhMQsIcRmZkSiNH6EDXS4c9xI7oB7JZYP/J3VDr8JIGMUvoBZ5X8Dg/RwgWt
+LmWjAd8JXN205PICt7ZkkPoKrBnc8gFyB7hwipPUIrR9RBEvEIOw/yM6pcApkdg
Ie+PFUYetnsWbBKhlvjCQPBGghVqt6pCvWkV5zxB6KJzw6fVXutiugZ2CGyADbFy
VY/bNCF3W4BlnqdTDEF9nA8hisdhlLtDOPXSGPuXH0xg8yKYl6WGaV4VvSpx4tth
qT5TJLFc/rLKSxS5EaEyD289OI9322UtS/N0Luc3mDs6O9uoSVZQrx4akiDSPuJa
VPLEwskVUJacDoac6Jto/SMB8rH96EFsx6Gbtj2DSzXRhKMVbkJhaylN2gZsndIc
SwRQWEX5Ex0q5N2G1FIl/HY6RFuPuUvc/IXpr+h9yq/jma9LdUyBMbkq7+n8CqTt
4G6F+Ulxcme7Am3aWVCvNU8R2xxxS0ary1SrzWsukHwdDcxP3hwfz7EcfDTXyvRc
t4V0UnaZIuLjZ1ILqnUE0kw8fbVivObJgV7A2TAL+MmWOPkCY7ILA7/EI5Fb1nOl
u9+SYABA0AL/xL/2XciIx8DMTdy2YgdCgimpoTt9GdEIsb+9U8Sm+0Sp4YtdSJMA
O0CPwDVdE15m1Z/9FO5tM5015FV/xguGmxyMS6N1syqu4mIx073WOnLuurOCw3Sb
77I/d+cgeJk2L+HmHvgAr+3gc9mfoukrRrTuKzjo/4OSFLukmgf5A49PWJnsklya
7QvmS3YvwPuipFtmvjA6QVBikrbzNCvqgWCrdqS26nGD8w6MdE+h6kioYYY3GofB
vClxZogdVIfzgwFMDVuI7d1XV2dm4X2hd8vMD1VvUkAPwD3Cj17veYUzyAZa1JN5
6U2be+Bp1x0Xt2Qkutm5JaG3X+OKRvOY/bn3q/86ZeB8EtJpIcAtNix8OTexRFZr
C7nX9ssRwojP76fvP0Y4oWD/yXFUqzB33S2fdfKI6+a8mpYdDtAn/IN6QG81JMDN
3Dvjm58j4uZ/qowx7sHgG0Sv7kQGJJ6cBajFh31a9pQjPLWQyatFp5y5I4UyUlc4
0782Uz6m4VnL6UOXOY19HKu7xdN6C5NLYrcrmQo6MNmef9HO+YPPixZwpwGTJZK4
p18BBUe5tLNts1tRfysudEMs33QsIh99x+F5J4jFjT+rrs4SAYi2H/a2JM7nibTH
xe+tNdSNVfKR2udki5wokgMpZQhQyX7DrZOg9Frn6lC2HEmLOphh11VTMQMDoLS7
Ad+n3KM5HbgXCqzyloVqafMZs71Jh0JVYGjyjgqpIqQm1E2cslV4r4fY0pAR3LXO
aFXe2Bl15U9zCUfK/WL7E9i8Lx/dpQusvukiS7c7VTzLzNhsr/2OpeEEtOgUKWAJ
tCcto7qQmOCvG+Ck+ugYTBU2U5sP90ACA4wp+LQzNq32pSgeXgsPevZ69fCNKfWM
Dg3xQHAcLNB8Jel1qN84YBSJPNu8gNjfeGwqhf6PlUrnaBt0FnMd1AKT4IsskDrc
45ZnhgEmuTMpxw3YpqD7fPLgcQbjfJqEtoK5jia5dknaZBhm1SfIJQJmRkxK0OdH
JxmQsXAVUWLeAOBSLdRQroUMxKxAw+6r155CrUDOprsP9ZHRauc4B3YnTYvloJi9
Z84TnY4wgZDDbEKzTeQxaNL3jwyp9uHQ6lK2L7wzkxlGxuDTgDt4BBZyLn+eS0r1
gAkoXmKkBYSXK/Gg89Qp2ZPLRV1i8YdOl4BQ/e5tF96+PaTQg02BDd8Aa29A0emm
iZ+zInOjXV7WFhm342g24tEJktamHFMSG0WJ9td0Gqv/z2wrP7MkD4VbZDFs49dz
Mq3V39vAoLWa25KolVNMGSAkAfMJy6Mr6Pd/MRbuE+INkRHrdPBEogK5/azznUNt
nXI3BAYUi93b5YDVXUR44m0E740deIJVYRNGZ6op3wATd+3uTlk5RZt1uOIRuoJ3
Y/XcNkG5bC+DPzn2MCgmxO4gziX5wGpCGjN2p879X+E/ryDPE8SxXdv/bRJtefRP
hqFZF+RXxG0Ea2xsR36cpI6RoQe8jqjkcRLbmBb4o/qsPZ8+BRkNKNr+b4H75SjK
mgtukOXvfv62beW24my5IN44BmUK+eGsAZPDmjwPljWl/DmglZm2/74Xmhqw+JHq
+TKxqPCHzfr3FCgZ0GiTMYP5GXCHkaanSY+mKEW5srIIxAbNLSNbF0nCXeGcmytA
qX2Lmg5ju0MWtU2u78phpg9UHZAeHlPmSPvMbSvXeJhacXviHpajNyxVB/SthEvZ
rCPYayVcXXAISqmBAwcIw+NOiwF7bDuN5OFfIqpa/5HAx8YZ8Z9rnYRJcOeaoxeZ
b7kkkrj5jsUqS518A7uPV2+W3HufnehK0Ddetl8jz92uzGiFcowhwwl2AQM3SmTu
RLp1v8lesRmKCun69WMRyzGT7hqe3fh4sk4HTYc4/zW6EInshPF+rBLJclkilWzQ
vmtZ7SPorUS+dBEgmVV69fms3n3T27eJYb0RyELkY3vPX4+S4wYU9bkD68Nf1pj8
lKzNC13MSAc9pqGbsJiWxFFjTwi0IpXu0nmtEFL4+kNBT82BX2D85JnqhqDKYRVv
oRxcvTcyc/aQkJMMlsA5uwdk9Z9ZS13tkoHabqEYNsMyS/RAvn0HxQtMe8Xvv5mu
MO/EXlE1EhwACuGoW0TkrTb1YcBKX26bW1IBMfQuEh/QdFLzZq4OgsxCv8Ky+P/u
9CYgE3DmSP3mpR2JxksM2V1UWU5Gc2JqM5ee6DjH3141TZdl2XGSKuvF6s5aZDAE
2k44+FIi4VeeLp+gfbHHB3qaed9PAO+l2LtfOc2EJzO8N2z+mxUgt6uQ0NlwjLP6
sS5KFa2tiv4EQJb4IE4gNXYkHexIEw3yuOVvBxWNgEZE4G+XsbxayJBENIER0BfE
JO2LL4Uv2SwmT+az0KmWS/ggJbKZfFEnIpqD0OWkvJ6iLNqPJKCwR0do7/0dSgjz
8vC/1ydtc/n50kOXSOjw2pbY2CIyt/FsND068b0vpQBBJWs3pwQFUNu6wAI3/g++
Hy4e9PwOg6tFu/1231r7TlSt7nh+EYUqNl6PGIoNs89orHF1jnlFlYzcBO9oM7UU
lzNdpf1ABN7XVte7h3Za7FlnedlXN4LfAe+jMSooeXLHgzscEcCWT26MBATnQm2F
Y2qxfOu2KM3e6AXqvvGO8pIcYSngG2JXujYXByaJTZ9+pPLp8m01TjQUN/wpXH3H
HtwbGJ9vQFqtgy1cOFfZOaOcP1zcXnH2gHDq0bhr31s8zM+E5SmG/GL6wg02y1pD
uW8dGVI5RaKdGf4PXnLqJTkBBUyR+EZLAgdaYgfq+1xnC531z3EMub2wvNIhgo2K
PQHd98+x/ojVY4lwst5+yfTus8BXtfZSFrCpUvhP5+iQA315cQXt/rSk6wotCaz+
kI9YExMPrwtfEp1leOfTSvT7/fbKvEYTC3CZXDVXd+LwSmmDcUJ+6YawOhwlxHlC
/tyDpysW9SzKJz0n9TWFpi5bqtBrqSCFIVjuCciXUvqLEWLcUwp8CjL/OIlSfWEu
nfqmiLnXFGxXmgLJubkM20LIEZIPMAhk+CS3R49nu7BaOQJeGV4mRkPcqcN+lm/S
rGILPJS1z0+osALPX/e/Wg9+lCq6C0/3X7/VZ9ow6Ht6Ihk0Ev8s/N9sK2IYfg8K
RT7HpgtdMq8+5mKuTCYIqkYedJia6dDOk/Gay8u5sPGjqRCumrUPcpE3FzjQyhpC
yXo1juAav1lE1LL97PYPn+Gpy3CC4T5wqtAINApm2BPgM7py/1oiwsokUv/Ya27U
A5cdriZ3MlppKHLGVCCDIZM34chnlMIZxmQN6HHzEXBkZZUfbBHxb8slcoXNrdhV
l3NdBxexATmN30am0asN8rTSsdypQ7rL5hb9yMSkisC8hsbvZmvet6goNrkyIUne
Ebj66ZF1YhhwZmgXT5jK24QmCiVJNJ1a680FnrZb7Igu70i/M8K02lz+q+kjuMHX
wpOLEys472OjD45Yp9EX7SJk5TCrxw/ZdmfnUVV4Wa0p5N6EMbZMauqEFVmkeQ1j
IFU9oF4qxSjttlR1C6Na5o0568oiNi9Ppcm7y6RdI9Mi4q2vVPWs6AFlcC68eJ7A
G14mMP73zJRCggszFdu6WfEGQtNyLEiS9yv1ULs1e7GzQRZqfLgoP7Jljam/6u4J
C5noNhqYG70+8cKqECxbEs9FDeEkjY7n3aFN3Sc/Zucwyh1XFikMDQ6oFIpFYkJP
mFCdkJtW32bM4vj79ZD/WYEd6+dMtVJXIxhh1+/2JEDxSnx0eGA9YgK2zuIZOgzJ
mMPpEi6db2nuEtuvANIMoN7Q95S3wUbikL0fFk9ee0EURm4eJa83WyHQTFDk3eml
vy1pGt50293zsZ8d13BzAGr0JvwMjvnR4B3ulERHnGmkk7zSJ+HYe7RsfEE4StA8
3qGeZDqYaxiAYdkKeMbxGmxjsOVVDjtu+KmeY9+V5/i1uCNRsrW5qGeJG+rcTWK8
PVzl67YgjZL81nWZe5SPYqhvfGL59dDE1OVyZ95Zu98Sjojcqr3SU5ILpOCrkCoD
o0cli1s+jl7nDI9q42quxnQ+7P/j/ETEE22WPfBFWPf6V0BqBtNILRegk3ECt1Eo
lKDBPnDEta8Ap0UxtQFEKteXT2Y+7pT/D5QXjo55nNHQy/02S5i+m7VQzV8J2BuO
c2oZAuuZ6fzhpIIUDM/4UdZoo5OJgszSU6CY4Hd49m4xdGX14tgHZ1b+2Y350Q4U
ZCi8+KchMW+Hv0TulJNJZ9LnufLVPuHtY9hdFK+Fto58YYj56JAEVN5PTS5mjhzX
Pn7LrHSfvkdLSCGQ7ZoGZMCybrtLyuzusfEVqZykHootpTStWqjaq5ZB1cYUbNeg
/qGUAWYknVVsOtovKoowv0hJfu8RUCH1FDWBA3flNsYisTob3lERRoxLaW0baH1v
UdI7JviReiUAbgIQPcG97gmC0jh9m+spdP+5fAfjCvUjRKwUSJe05q9UsPWzFeV4
R4vLhcEG7nU1rld1snTBAFaa3+vRYu4p2xA7ElHS9QjjH/NA59o9I00tMhaPTqYg
4RFk5K28l/gVYmNQuxdMg1bBarb975z3QGuUUb2WIo8MUCPrAPGPRI1WPSk0vjC2
x+cYOWssKNw5XqePvzUuGB52aMLVVlGbPy21QtHq08OlSti9j/6Y1yXkBI0+sgVL
ryrTsf25Qej52uSy447YMOHZYrIoaOxz3sYh7oqA4mKLv+FpaJCXXRQZXZnzUl8D
YTbCyRZPXEt8yCoQkGw46otGKaFLPOFCJf9Yi+jg1gqed8s2aLbFD4aeQHZAc25p
chdd6hvlNh8oVgb8wIlAje0jyvy/IS0Mj8cT3lhMBp4S75L6euuXn9jOZ74hnPKS
+qZsA4QxYVsDrfm+cA32TKNoUGbUG/7kHujBIPd48UW9ql/LnQbDziLOJ9sGsi2B
hVImVYdxqtRd/E5YrcoRHMvdi7fE603xTtdhM4lpUhXqJ201PNVSrPUeIZEacu2g
+/xt2xcRWthgUYZIb0w3FYyx7GH1EkPgu6Y9QP52lDClcIBpFx7oDAZ1VSqmUg8w
BiViaU72DhVMNAWJLHdz49d7myViVG1E5UCNZXNTV0xIFJd3h7miWDaLvNYQ8jy6
tD/WuvLJ9LgUKicgh0XRaORiEhtB7m3N19r8BWReqPa124XWmjfNHQnXFUKVrfkL
JNuQ+wG+nOl7PUoklhXIime+x8VhFnoVE0ttdwYa+zq17umL/t94hozNoxdxpEuL
NuB+MymuSI8oyKwxz3KnRuOfd8cBPfTlm9iFnU+UqH5b62MbY0tcZpLdgsw5vTvB
BNdzZI8oiRlIM88xadcJfyEJBBvq9rMWcds5DLjIuBmPusb9Ogtqq2RYCRWlOPkB
uICQ5OLNAZx6a7mXlwJE5bt1Y29DWoC4Rfq7gCS6LY1Pg5dNbgyh1tuFAkQPz1vN
MEdfDIluGzVjiE5vfdIqrhyxXngHyzbhUXJj2TUf5jNjicblESulbDrPQ1H6oSna
VE6O7uqxTmIaCCS2RzXfD2u3LUVLyBwrW6JpmCOeQiR3FucUX1YarDzUVQVHtERX
D60GMNvKkiM8rfZUwa8flXFxp96Ec8fkX4vlSoLWzbLkZxnuykr0icjMU6wInUjB
Lq6xtcGdY1TixiO+ONxZ29BR2lNIpOa4qgr4CVOBU77mM7UewgN31/+t8kUSXM1p
59BNMT2C8rxxz0XXAOXKebMMj4jgViculXjd3l0n0z6RTIDFz9rYQ2e216bZw7f2
gPeWvBPZQ+JADSHs9IcAAtO7ZgYucnQqtpuqLM66O+qOu3ieW5wtqG3kam4CCgUn
YfXzLAyiTHXJMaybsDSueA9LEZ01FcBdeU3WfkaFDG1N6cAgzlj1OQ3sUw6ncHJk
f6SJ7lmAZOwb9+/xs7odrqut7wygMT7S2UJQaIeYaJ2IXgH5eGu5OrXHgSPt2384
PmhyE9CtS0cv3NIqxG44p+/s6kIpem/o0uNUBOxIEO/X3a5OXcozBBi8zaOXzX3T
8H9jhIfpfJ75t5AnkBumJgJdSIFEMxWGVEIPaNtWeqhIBzWT9UhcoAmD4TDNKSQ+
x75u9eXGjlcF6ZlR6SAnuRNlUXfZgx6EW7z5aCZmF0ax9uoWKcrDuE36grM7hAsF
dZ4tDrNcf+bk8QmcM5Oq1pWBNWLePxRbZu7/wIgZA4+U075UjvraGQVOxDBuCxof
AJNSmiGTFM8dzPAYmiJ5ecKkJuIILk1lmd7+oJFp/RnVW6ZA3GhZHUSz3MXqikyL
O5jjhS43Inzyof5U6KM9uon8vMzyZNVZfDE8Rec24msYxI+GfxK25s3Z6xr42Zxs
n0yRKrq3XjGK/BGHQxXpIH10r9YF544gjr0DN2c8q5Ud7LLnm5nCyKpzJr7unl1G
wDsZcmEeeXzXPYpNA2nOeig8mfNVXcmodiM87lCnBJXlDjCyGgdYN1MDfevHUi6f
RYwQoX564LRyS0zZhYtCZTFSHJQyzUM+GLxrM+hT/066XeGjVSTIK3hkmBwn1cgk
djQYtXtxY0Y+nZeMr7VgUJLcXSAucX71EYsvA7lWZR4s8W0rJM0rndy2Y9MAEkYs
avNOlaDuFBt9saIgKzCpwvHr6KlrS9CjfD1Ma2B4yXSAYwEUB2o1gtR1uUCuIlAc
4L+8/3gLoZM4mUNlrt7Vn3cb6YcIgQGnC4G34KEo0TjQMNfXGIHsupnE32hV+W4a
G8XJKLvHtrECxEhqWqMFp9KYowcUjmslLabnwZr0OwH7egXs7aQq95FNBD2/Kwu7
GzBLbHcxOSbiy9iHHM6AQJ8o0U7UnHJAm7xARFB8ImAvDHIfR60UUzNNb3cnqBnU
GlrzexGlecmuwrHh3isWrLdkqdSS4FqvkjkMqgYGlrOXL1OjKzLfsbNfV6blM52B
5kclkfj9sQCMwO6wds37YSr0zHsgiWmHZ1Er09bGPNT2S/h0+5LyuRXYDmIAydmf
0gB/5tMGkW23K8JGX7FzewTOd+rV7soLUW0w7XIvkYwrOeJFoTryCul5Zto23SIi
wCy4Y27UYKv/zdTw0n+4b3k6Urn9QSCxIgtJG3xpRtGNc9ob+Wzz+cr/YDWs6NAp
b1rMBtC3UeCnEw7djB++ojSwLlk1U+y/E1UXXADzCdJwtXK2bSTRNR72Mo009Hi/
WYbPQKG/Nt/OOIHNfY6SbiD3HSUDCcdrcW2HBcYf6cj9qhJf4lQBmw9XvH6/EG7G
f3gGaMwHVJKRBT32B3Dn9JQ58047hhKibcytoMb1/Tfcrg6XN4jlmmJ5DNYMc1To
a6dq/spTsNiGlqDjOkaKyN/gvieddmGhuWYfiGxoPbaHV6Ws5AX3C8Zty7Ld9D4N
IdgLJoXgkKQbdcqRImNofsGDikNJIuPhzg28RAQ7CCrmIbrnuHgDpQehK0s4bmk6
BowTsv5vUBliyKqCiinlzkdQ4L61C77//1aIDM1khM3f6Ts1CH2S/11PmPZeIzVU
Tq9Sxc7qw7XLMF960RPb93Q28NxfA5BK5Pq0d4LYcIjmrDHFeKikss4F+hx5SNI8
NEAOWsQyNz0ABC6xCXoF1I9gwr5YpZWCxCM2wmKyh9TJZ6XfmPCSglz9OB6Nrg0o
kDR7/lNksuYdcmSwiq6JCpFzzE3/ywVo8V/ThPPEblUPz6eJK/F1wH5v0YG/uY5l
UpXGugn58j5p9Ej86jAFQkrT6oMH6upr76eEm5YFKd8k2Mdd2/DX4zbVHUZjn6r5
0mgOuGqCkisQX7kXPZFWpu4huhkxis0ZSi3cBdnTNq1k47v9NI37sLbJIUURJpjR
i4PFjam3BC/h/ojPUSCpNcMPoOA299fLEtrQlS24afJwEZ2WPJNqSnzY7AEgdceK
PtRyUKjKK9rQKPPoEtBlWjoAdL15cxnj6VJ6j8eFUuNqbfhSBgHYTlh91TGMpWg8
FQYtVgND4KTgsnV4PGuDvuD289Frjo5cTBJDQO/H+VJ5vra9PXpjlfoz5tvguLu3
3KvDi+jHbGMUzkM/7aLU2wEwHwybgvMKrFWXbhheEEk+9+MKwIOdNUhaqdOEELWj
fkZigSI4xzfHwVHSqfu2lFkkT37RurpS4vr0wz1CiID234VV22WVD6lYCNz6lt6f
DCSKkHngiXWH5iD3y3GXBAm//I5YOlXr+lfD5znjoYjt/Zs1fjAf6wAshQFJAYyE
VOuPB/osSKPm11HjP6fQdFbbqJdQ1dI+Z5Ab9EY1rVEp4QWSl04PC2zEy4wwF1PZ
KiFwkx+W9838Hecf5aBBOpRIvQtAtVdFx9iNMoooAj8B19LbvFpe9T9mEdEA4bz5
cuRyMKYCeOVETEhw4Agtbdpe2YDzNUHTtRc7I2l8zokqlUv9EOLI54WJRygFv65l
cgoYLbziiZjqzcT9qk1kQQRzgsNHvPSs69ngH2zx/zbHNp5Qz+FRztJTVUYwqCz7
lurbwqwnLhrRRuLu1hysvEa+bfuZg/WYhVc+DUJ+5/ztZczSv/00PS9rNRQe6V9/
q/3VfZVWu7hwZAYlXrTdplLyS/xt9XbU1dkrspLlWmZwDpA1FN/OMDtKyxoRjk8H
8Y6UC2a77ARueHVJAlHEA7UEX8hbJxxi+6sifVfU6JzPO3pKfgAnrZvm0qFhjQgC
LSdujUZ8S2ATq38ui0qtCkC7NtyTGQiySa2aflmzb9ZrJOpDm89LJwP2Jz82J97M
DxbS2cXI5xuGxx8UmUEmzWoJp7qKIU/q4XHxf9WIgeXAsXbrAPj/GzmLNuuBLuvy
EFwpQRK6j9YFAvQbAT+5GNOhmBGDL/G1RrGrqinMm/4rpklGD5DuX+qZfXxEHK10
B7GWNONoR+a4XSQUH+i/cgK5cMcw2XPtHYiyzrkP0LP4QW/O425byxqU5RKkmLAM
I3WVvPShHhaAwYquP9rstUdsFscoMHaC+pc4TXLKFget3EjMMJYFDKD0/fcvwoxD
IGt1x90pCBljdwicG7m4zrUBTtJeKYfHbuDJyNpkX7+T/nZFOqxtIepSAeDtlfc0
WZArYh0e1YO0OA3S5tb3bV/KPvg06Ynl0cIL6TH8Ik5uCgIL6hs/q0LAvGugTIb8
6a5o3x8xMsrCD4Ow84cPjjLUg7yYP+ajqXV/6otmCIk86frvuIl4VZFQuT+PoFNO
H5OgG3M5HW+50eERDV7MpoTW3rLxpA8hGb9j/2eoqstU0/5qDxQXnfoq3ImFRShb
KuiTkhzhUWtRD5lmBbAWX8toZDiH6OFjWL+v+qOvF0VqsOLFoSo8LDf9Suy6DNXB
vDGThFxtCFXHDSor5GVjclCIYIeN5swmluV02LrHXYgQGtnT0MklDnLdD/7UBmDk
Ec2Rusaf0JPs++d6v2BIjGMeiftuShIctcP+yC8k32gKNHnCeNCmmLwZUjWaoJe0
GxP/ZW5CVCnqX/LkRK19yq6fo0iK+Y1mB+sSUDpDi1qQSHUYY6yYATwemYvnoRJs
Tt5Z88hU5/0yKms3gB/uqFvs35eGw5vyLc7InrY9CKfAbu4FJOL02xpdqz8YXXAW
YMKzaFw8ZBk8V3vtuNCOPBV8ZdZAGNMhhLDlF8OhNT31zB3jDn/8oLwazavmzscM
xIxzO08sipLjXFXuYB/70GRyUcPqqc2OD/IF8iXw6NF8YB+VMKE/9LdLLVqo0UXP
MoIi3RnxxsSnTZXSHyIfgOZR2LIpu1+oLIPz56GtUDw8dYQdp/EeQu9gojpb+BBx
ihKPHPWgVeAyotIYbnT6za+/ij8NJnWAtOKnN2a0QUWAolsPocKqHX/YbQdpGtEg
dcDB1YeL/2wcltwOELsOmHMgZwwFSJKbK2x8WiQfP3sFNdxoQ4op9gl3Po6/g4kD
o4HnjtzSc5SSLdwUg3VAE7Oh6ZQVqvAneAo6I1ZPYMj+/EVcKlKfVi5QlFgmw+Ob
2wyeJffRiCpIHdfHmRtvHwvPgZPq+kyfCnE4NwR09iACzmKuxsB3cCuLxXUeRKRy
6yjS9W2DuQCMjdJW++dxxisYLpnpb3JIxMQb+40/XfH2edC7j+h6fF/oC3mPxg/c
ksUMn2N++HHuhHNByVKdUfYywx0IYeCZdF0IOVn3+nB1OyWhgEI3VWlbJvX0GKCz
VdA52Sph4NOKNMtdrAGF2holwhPARCk6unShNGRmlx975TtBO/099ygm756Brx92
6s43CKnjHqmTt6GspIc/XR4Bpr64oa2ttkI5eKc59W/lH87NlMB90JiQIbTMCeCF
CDiXVm8xTz/r9sGKUwulF51fFVAeq07o0sv0XVIO6w4jCm14Ne1MUKd84Dv6kcv7
4XiDvPcigmK2ZmOlThO1wwMcmCebTVdbrxW3WwaVCYzlkkas4g9NSjsNgldj68B/
RoDfBroE72ydMfT32ep0ESk4y0Df64IKsLWKGq5qTS63BX4yp1W0vn6DKDcc9P1p
XZ/h7fthC6AVa0aTph4nVrwwhoao9Jw64s2wtCRR5NAUoYaYgTbS06KJjcwp9Eg/
Mm+ExBnqQP4JiYZrL7xUfdkoVAs5o7lMSIsukAD12kiW9ryn4TF3/UGs+fNigDyS
bp+DEaPeJiVnkKMI3x99ix1pCcgePuAtBbSzR5lLnOsf0Pilhd33BcH3yJCreBUt
KaBEwM6QPJ82N33p4XNp4FP8OhNVlu7k5bFU5/TSixoxtbipHspcElALfL1WSp8E
6P3igpJFxd5yRUBVnGC0Zz0HQbNbV0QbUVpjj8wy0YxGhokpYwsp3BjJszn6Emg8
3Q0eHbGyE4JjllaMahNhlhlB8wNGMbYMDGYefpVPwpQLpv0PnxrX74vVfarBvKgM
qqlEDHF/Gutf5yL3GHlCPuu/hyFeohaTXBD9ubyAV9clztzFr2+YfQoeGERQM5+d
30lEkhoYsAgNsYdpffqY0hSMtMCiTifrEPxsPkyhWZq4vGQ7lNDF1CNa2R+U3lbx
VlpKNKO9DduAslKiT/mPVpr9DLfFjJLgAgYZhQNeCxBYlGaY/qZqpbc6c794F4Rl
JWI5XutRdoPFJjh/a4iaytSaJIUI4TBrnOo1/NEkIBuBCGdZ43Gbdo6pGJ9dPVyQ
ybD9+UzPc2TsUt82FsoC63QaVT5EsjHXfQheqiBuDYWFHu9/v6KoxMMkYvAX4mz5
+IyXYrplVcA8ZpMlZRbSABIrw3VNRQ7ydFA3qrFe/ckRjcLRSCU9QCux5FONFzyn
ibz7ZyeVQxohvaxdg/lVD4de6DDXQm8BaKDJ3nyQK+kGxL9K/W720NddxBjz+oS7
lYJQUgDPk1pqCD3MSj2gKEeonX1aWUxa2gw9w6MTsJYtL1neKyBDO8AMJoqf5/5m
2clEBw9/QYNRwXFOLRsCkRQADjxwYnbKpeEjtUZzgwpxi/Op4YjadCtaftpC0q14
ZjGY4i7+CHsHg6vKCvcwP8j8y1fUjMqDmVNpiiAjUXBZ+QhY5bHAMdvck3Ie4aDM
C2pMQDR6gsj7fdtd4Wckagm7cJrtQ2ojuOQkUEzC24oRsSfL926flO3ia8W9rzJh
i6PhKohw8PHEVUTZF9VncxcHwmeW4584pHP1V+sl3+IxHwsd8VEzyMoHPUGGdKlJ
mFd5v2Nc6eOQR80f+T1D8rw2Zoqbc0etRR2OHlUww6Tjl3IsAZ8gczzSUi00z710
EgmBV/DZy6OTYDE4WcgwE/bCuTWbk/BFCJ0B4miBnjRaVR0b4wudwZsZny775VW/
INwu/orMIWpgdHAMDHkIYp9xXhHWTEbpJfmlDwjsUSOhgxsSJinRCoHJitEbCqbf
h+B6qjrrG8G1ZzBxoCkhdlPAoNC6iT9viXPFAMPI/C+ow59u17lq7+Q+WMee4Yss
oY9X44lS2HA6C6yNcOA7AXO1oox39djW5KpwhxACgGf+3X40LSvSjPmQi3SJajU0
UW8S6Y8atxdfWOS+lhS2Qx7pL7OCi+KvqWdb19pT1fPq0RIfvzWWDFInOLicedBk
YEWu91I9Ls0cMjKLjtyU27B6ndLVk3JXiquPE+hFSJ7q8jjOgPDWv5BPZgRW4Ngz
AaDPxGor2rcxGk+/1+6PPjtokvwd2UqrdlaxipUwO0Ns5xlX9diOyb0wcr2j0+kO
qj49acu1MQAtp1HIIY723/S7tc9K3odjzR3fJx6RHfKXIGo3XWDykDJTLkxgCcnq
aHn0zG2V7qbRa4wKU67s0nhnTYqiDsiItnp5Z0QWGccV+utkQNlsOwfigyhSxrXq
AZV5qPiGXEfc7LguT4Pd/9I4R/uxeg5VCsR9SWekI1Q4yH5hhTvO0mUmHAkDaZ2J
hcaXVHNNNYrClsaEZX2eY2D5OCCZOhdBYzaO0xt79Q4j5/ccKOfMY8kfSWz4eMvk
e+v6yTC5U2qrseL+bCQh6L0ajFR0cxiH9wG4QHwjjd8GF6IouXoQDdoojXpfvY9F
0Bq55EdvrczWSMhg2vthWn262MT39M+wajBhoGUCHYfpX9YRdmgbMe/K8vduRNHq
do1sekNxHJ/5DUwErftSfkivOEprOFH6lAQbl7t0YGeSxHgtEWR4lyiCT2SB5/EN
/uYAgkqdQ1cdjIH1r2rRCkT2PRD+GpoFA0sfIZm0eUvmLBAgnB/ib58bmbzbKoN1
2nTZ76dpQ2Up7Pg2wsFYRZBZ7mPX7UzJ+U9w8UL8AhEt1KdknCK4p8g+fEdzv2a3
GmxO65qtk+asrlXcJatYzv7l3yxXu5FT2pxB2ET5w3azA41Kj71pcYhYHYoi7RFR
sANIXQ8l6uemyyxnGEOteDnIbkV/c2UcaLHXe9Q4sv+romRczOfmIXT5qpfS/aB2
YiucwDznd3EILPAMowqh6z1mLNrUmXNvZaap9cJ8+55glrkh9Oeqb8jL2Hj2sCOa
tPHoNoBNuaMsqvQy7Z4bKfN/tclpiB0wz226kdJIhH1DOIpWNJHCZlz8Qks0hqZ4
19ugjei6f1Ihj0NZrlyWKJLFvHT0M3AhGsUyiLneoQSiSXRX9Yuq0H3F95FcquWJ
2thGPZA+bxJuzVyT1Bjt/F5ovKStGmaBcJ3gWz2yLDFMUAa8dd8VTw6oN9G3ij2D
AufQn3a0cZEa4EVPP15a1En38iNgLaerFH+L0HBoJ8MSBGHkhGEJMvEaxlrtbA30
sOqeJ0RjjYrbZUkG1dS1sJbq2AceoXish7HCIuVYkTTOrbhfMD2dskagyKpdx7mN
dcxnLtYFR2YRtBqFgkdGf+CeuIYUcQqT3JOJIRlEge1MjEiTKpxpVRfLdMMQjshQ
naA51mzT5Pv927G6CMDo3aWr0B4iJl8/36+n/J4TGeZrGsB31bqI7ccqCz7zHiXV
y3G2yXbJyAGGLC9EcItBkaZnXTiEQw29YHvQoUe4Y3XW9rcvA6Ctc4ReV9FPfTCP
GdA/8JGJi7P8J2u3Dc5RDg5L/fNMovWmknAkbyherWRPVjJVwpXW5Sd2VFxsGo0N
xptpXDTgzub7Ty2xGUi9rU85Tb+Ja7+syFwgJyxGCAAIQMZJGPEMcyEmwrGTZsmZ
p4iD5peRZkyuO+Xvaro376UZJgB9EYp99HVGBZiVJzuOi9cOiu7vaMXcgyV2RGwL
iTWVaq77jibQdy+8aGRzOByK4/k55oVSazalC+8eE+PlteI3+MGK2SC2/uusM6QZ
AP5lz7eQYMi/h2V4YycSL0kHat9A+aKMh0z5xarmGes8H+PmXjlYYNraFO2UjW2E
4YClEZ/opUrNXy08W+YxtTmWpeyH+Dw369NxX9uGf/UXH3g3UPKeLFjxZ+5CSMyg
9f8Wv88Y6SU6dkVRwEOPdY535grSNPhrzCnLlQs6b38V0dsTReZaqT2IWFSxH9dM
BH2eEnR0cCJfvSXKZW4u73r98WCtD9fcuiBom6NH0bQ/odmD/wWepgn9/eWVL1tX
yln+U2wYzakgRFDag+fO0b/7bqlENkBn7YnrFyL5hH6PXVvuC971y0MFrx63SgI8
t6Sxxo4aerepN3LO+R85kxGZSl5qtXQpoOBaMNVuTAkY7D4GeSCj5bylQ09UltQN
xlHEp7Qyr9s/JrdnQ6UQ/IbcIOHPukWkn4VM+aUeygL6z11j5HLm8Y1lI1eVH3QZ
I+oY6nHf7TZFKmoIVJbpLyLkM87hBOuAAR0mj5SP7lVNklY3vqLin77/VXNkfFUY
4xEopJDXTuaMbb5To0CxJd31ypEixwOwBxSErZB7bNZbAYfT65oTkRiDLp60h65K
5cjxVgcvDR7d+vCCx4KssNsspGsjQocPP7RrzDgFNLElWZrTNc/PKGi/Pli7XU/i
WWC8SPv8MnQFGKAP2BI/GdWXW84oNWDaKTiaAhKgxrU/R7hZBiLNnIy04W1Wgyfs
FCu5TkL5UziadITUpXz92Zm3kKyhijPpFRXrVwWiO+RaYVpeqgo6eA7eEpLHOnxB
a/1NMm2Wl/8gImTlIM8ZOh9etgAhJD94wK2a9xWE1Qbi82C0xHJKKKFth8OQxW+R
XGcVIV14O1+rrNFD/URTpjSn5VPKRxpXnTYxiwj7UbcEeI23svaPWVsuFa+5nwO9
Rvutl1tmdfdc7AOWYvnk/vd3ZFTFqEjbbXD0WUXbMHgYJ11ZwzgGMtUcZNsKExVV
2D2DfTLtYCqvvFPblDDWEIuJxRGAjN6csAffzGR97xqpbkKSdfE36LRqOxx3znko
sN9zk5+CRbdAJtV0mdEKAh1SFRT0hqvXFgCcj/g70OkvSQ81Y1dkrAo0OKLmB0Xv
IbrD3iwL0YctSycWpOSNVYC9qfnePdxWEFB0AY5EljJrY6+k/drrt7Vz6ZNRB2NH
hNTCbU5MFBgdvWaG0eAXMAUFwfwYPd2AJN0GZ08kIWpE9h+AK0a15gPkpMltTdmn
AzJ68RBuDp2XKrPJDENVRAMVYahWIO9VwPl73x1ELlwQHzqMBrOus+3+2FheTpzr
GhaABGyYQobv9wHlMCNYww4t+q8B7Try9vMn/iLg82zzFiTQCEAVGJCzo+8THrsG
ddhg1xh4YlydoD2YApAyHCToGt303sEPeyCrO+/E4vDRld/9ucc7ceU2u0PHB1Tb
dbw0DM+KYLTR+BvkI+MNCowz3THoBTqkpQDa4hM/2B8PWx2JblFaxZuRxZpOFcc2
VP9ouzu/TGUo7IV+7NsLm+o6s366KOnyryPKyrPlEcRyLPfE8wVuJaJxCQKW3ikH
VYXcJuBRmq8fbqxFdSYnUUNnMbyrcGsS4QnOusdp0LLC+/8klbcCRRMW843FXEzr
jjOYOMF/B48TTI77sRYdPNpIbQ2ZOS/W7AFLGZPjUpZ/dhfCs4UZ78iBzFjnyfA8
Ff329B07wPbdhLbumvFo7+62xWxcQRVaz6Ll5PEII3i4/eeHjkjQ+GZ73rzp4zbD
sPlgpiYfOOE7xowW3jfH6JGfsA8jX2xLrfJ0/5m9hkOp7Oae8fVCT+ndp5/vibqr
cncFZ9iZTp6ouQr3G1blkXF80Key1TrK1XY4LEWqwFc2pSlq2HydO7iR8DhXuHdq
4j6SS295MJ6kt0Ftk4OkwhiEBiysONAQD0zAgG5H3aqGNf24Rr7ZpWaB5AaGP3E5
jp8jcFLEupSIIRwKMJ80h26UkL8YacAUUg50oWgA33GWMr8BsP86D3IPAr/CQVna
i9o7V2y73i7BZgcE1N6lwwbt2SMh4Vz0zohe7AE/xeb8g+19BVs6NiOqeqF8oi45
icwwJaRv9rsH5JDJAi5a+FbnzoayabBgP0+u2MQ+0psc5QueY0pK6iA6+zSlfEiK
kVa00Gt+1if9Ay30c1oqGhQpw7rzfIWj1iKJr3GFXSZgeGzR/+OhOl/4OI5Vas9q
PsQ5vD8Q98NV70oxzojks9FPY4yBihCdrh+SFubqkik91fEhd6yJaaMDfEfT2xzl
IcuihkOHrakMKeeBFl+QPOVd/kf54pja0chQhASYk7EEzd8JhfYbcodzBWfHJQu/
hlYqy8Oqh/9iKDT32kUCZY/lNyqVcKBBxBO+c/TAVodPgS/Bbt3A1OM8cPtcB1ev
rIAAt6wwmI9YPfE9y2eB73n8z0czd7Sy7gXWpggmjzucJOKKRVVwTqk8pqpTNIjE
MAMf8m4XPEmbb5NIm+4cLfYQv8cqeovkNdTGls6hG1vHD4UWTkG357JTlPx4MtcM
EQhnynV8efd/hFCjGBc9ToMFxbN40dvnW00c3CSUR//TmvsNlyq8GP/kY72y1E9q
BNbB1APM4T/A2aUWBODNJOoqe6irM470a4cusMNu2Q93dKRlqqJmeGY7spkYZL18
5Q83gHMklhKJtizeYl4xS7ZgyE9UyG1aB4YgCSU3iTmU1mKPmuIdAh1uWMv5Xymq
V3u51crSwS05f9AktACjOnEkciAq6fGk0T4dxm0o1o4VIhJqRgnG5K6Awy2CnQqn
9B5b3oxWJsELa2ou3L6dC5dUdyPI0gx7cqDK2bY7oPWkjGoNNcJszMTEuGpCRI9g
V98dxXTkgWbW9XpajfPUS89WFZ27aBrtJ41BF7hyJqajdkHzLx2leToSidGo5Qmo
cNUXmEuBD4DNz6AaubCWcY0qobhjMTpTz9SM4qE16s3kxbBWga27DVH/K+9AOlaQ
gkpHRATwqfatt2nlUceaJA8HpUO2UQdgruM1llNl0B8oX4SeX3LS8z4tUg1CiHme
eQWgcDtrovadpb6MzPn9hxjedTCSSoD+JqF7QiUF08VmdA+Q6P26Jdplrj3T6XKS
dh5EK0S4ckoOXWFIz2vZBSHgvmQvTv4ErBEFM1eQs3lv4RMBxXocnYlCLvlITo5B
pF3ryUrSDc7oHPuShlWDwYiaASCJZ81fbrpfrgtWDHaTjlpK1oy5UCRSSMysxNzs
Pk/BbmVuffpGxeyWJWN5YCoLg+9aucRFPobTeTpkmVphIDbrAi/dl/QsS5u6mAN/
9vuH3GwqvU4BWh27TPdR3UYzSG8K37Sv63StXxzTB2e6sBDtT7dZjHj1jfVdE1kG
D1xvl9pIom0NH561JTbXq1mnjRq3EEUOwZN47vuNV+x6OEafOTh2EaWcaa4Vvshi
ZoEfGYG9mxsP/+RqfuugroDNq3p4gnre9MPWzXonHnOxizKDY6QOWUPIFcBa5SSh
sPlyv9cqD+NK3a375tXU7u2036hnRP0277RQrgO4aXg7PASJiGevXjUeQpqNPGOm
HeRCDORV5c6JRfhHC/6OszdpsHIUANiZff12M5DuQ7zrPUV43jZWPveDJckUK5fu
kSJwdHAfivXrung9w1CiZhsiiS0Xk8dQWy5aJWElpT/EsioNaitQXCI0HKlfDBNg
u6d7nCWAVRfTfPkePRCOtZr43clk3oHatLs3pk4L7wlngfc9ca9BY0qzBJS8dvbt
SPYynnWFLHI6J5jGa/tDdTIIi+C2XCXXyioCnZw03gIwiHyul5I4n9+RqJK3BCGC
RadsUp96/1vLyphjtyM70+Uss4VJKr74MAyLb5fMkIXMkIixWIJ/T9dR0hM8f0dp
czA/cnwacVmAgYqL7R2AGGF2wAXCRogftr7k8ugZdZNWGQSvS84fdJKityojvXRC
VouPlPOv/OAoZbqObxGHooaMmAEUd2dG7jXCwN2Mwg1fg9cKM9/aZL33N/maKUm6
hBTct84mcf8MZsIoAKAt8dBSvaQMt1i79az/1+WKwwGxxrWlGEIs2QOXpxwTkMTa
cg6XMP3CzXFKCqOTyW0OkmB3WqF1K3CIME7S0p4SdSwAm0nYAzPKn5PQPxD5eZeS
AIoBdlYyzeks/vyzE8lTnZFl2pIjanjN/ILgMUSGTI7jpPrXS1gZU+XUOgqxbAEH
h1kacXV+hQhoLmQr/MWS7GGPIJj8yIKGTHYiEAxULTn4V4ISIr4nFsz5ajz2VOyU
QCMiqzjlHlzm4N6iFJWIVV4qHG8MXoRFNbNIz6ASNvKQ/enWo4dIj3pu6zvVJQzQ
wt5gw3Y7G7xvEXMZl0Fi31zpN7AM2lNTnGv8oyz7TvMc9shlJWvK6Aw/LbnNAppA
GODc2Cn2wpWSYNVmSbxKg9dW/d0y4BKbeOiLMLbUYuSx3JzbZ8oEDHYAY3IwFMRH
BcFjTBumTVPyZIYXAVzHZJClEjLaOWFhMdW//IDLvDnLmTybPE/Z4IC/O7ammf8n
kPerxSM7YHgI5L9iTUo9rbNaawzBFFzgsG3kAfythsh9rp3iWeQ1caXDoTmXtDe9
2v677Dg31wMOqIAi2EZYi2v5TIafOo60WyHnouVxLG010mRl3ixU2u78Xd5TVpeI
Ndgw7c0lQEMT3C1ea2ynQ0zf46KhjMciDkrP700QzBaEajhOzMfS4YDeaH2CkG/e
NiONQDYQUA7F1D6+yLnQjRpYRZV7Hbjndo60FgEquakAqKLCC/mx1MW57zddFcv3
JCWEdaOb2ZwIe6RmPJH1hh89aTcLXL7KbaQkSbxeTHx1hKY//31adllJtaaz4urC
sFfNE+I1d/vXO+IwsS1t7YVwieWC8ALt/JXH1uXBwosojgWOc01zuexvU1rvTSnv
QRJEhR5hzRV45GLJec+nDQm5Lzaijka6A1DT7aLE5sAjGC0iicscNTAkYEsRNV3h
4D5mokmKkSL64VVPr/It8LHufXyy+NbCPLvatniqQs0JfvzkHqPUGjZduxK2Bhk3
uHRDhsa/LoQFVxla/U47CglPLNAW0gYMskd0N27uktk9dM8e6QIESG2ZnerlnWdx
FCWUhrjbuZ5tg5XJtm2LPM1Wnc5RKTc6SQazzp3F3ni3WTzz0W4iiVlq6Euc7dhV
9ii4a7GVRg1QYU7EswyM+RGUXRSStS7szEfMeCQbJz+zE4ueT0s8xF6H0Mw/l5lX
fTWVA/drZZQaL3baOMyizn4ltTS1DbHUPghYRuYso55RWJ8I6urXqG72yhm0xefS
IJzzSehzbFoE5pSO6E+ezBt60qx875os7eWKMH3vhoG1wg+yYvZlD3OHGg8LfBPi
DBYQzGGsqZjzn4iDWRKegYSmAhqRhYvRIUxcl4T6i15kNWO9okr3EAMhjynFqzeL
NmICYWFyb6CqUklaPmlkg9IgjJuvlVNFiKvMsCyEwIyR/WT3UU3isycbwiQkZgu1
tE/iPCW+yDOEyYYAJqQBEIg1MmGKZ+BizooamSXCNidcx7FErqmaaiPzXo0JzUGR
GpkfGOysG2s1GOOlIaQdOMrs3xutM9vDxkr/ytEwaN3sWKBYrYLuMzHNoCbbtKqC
hZWgK+N/Cr/t5Cl7ZXy/Qb4QWS9qC+MSMO+r+jJZ0UwF0HYoSdGpHGGxEsQOWTpL
z5KdatcN4HpOgc7VYSxXBW036o6kHxfzWo/NexKhN1BG6Yk8D46h3hxK3YzanpEq
dCx7IFA3HecYrk8KEZPk+rwQEZYsf+iJ0/xPexgm+HYMG1NYwYMBsqP9glAtygD/
dVcYnOU3kr0kT22yV6vcxMJYlbK2IV/yhcHx0O4SjDeTLY9HoKTIQ7icATPKm1YP
YodLMfseZDB1UwyJWcMnkn7zwRA/QMKOcRWFkFSnFSNze+CtxxPf+n2rIZRFZZVS
v8vpN1PFubMEHUy9pxwBtfIcrlW7JXoRGB9rZXBNz6IYyVZEJj1yOW8Seew69YbU
ox++AfcwLAEO2wuZIbgETciKlr+yFNCKm7K36HR60tU4owzetrqRq+H60CObF90w
qTUS7+m7bZ6cHJe/B0wF9zqSZuPFQCGejfhDZqSJskYkJwsAnGTVv2P0kExqs/u4
lQBkss+q/aHKYHiZ6dFZ62mU1Q/YLanvMjnnNUzs/+HuetRE3N39tfWJwpOlAhyq
o66xJ7LhgMxb3h8uK4iV1QQoLqkpqcpNBcX+ec1zstCPs4dDmwlYcJDNgaYpwER8
CHUd+mAfr2XJPMKivEXPyWZRUPiMv4BupqiEBY6UAn94/z9w03IEkYj8mMtReOVO
3YO+lMQ9uQHxrk9IIf6HFERDLCo3KlrTEL0BtvwzDmDBoHFfb6kUGIuJt/u+sCOB
YiNN/ynR03oJhxtnwrEpuWsu83ZWxdCh4A+0zLahp2uRl9jrIIek/5mGWBe9nst0
3NaPUf8xPlyHAxbw74U+P4LNvWGiYkRSvCoEZ5tF+MG0dBI84YIPMf7WESEbJk8F
9Nmr5dmNFyFOZ2j2ddzRobUfOquE4CTGxjQMRHbOyOJC2nQrj8XgP7sBcPVOP2fu
RqaqQwaIzfqYCR75iaGLo9E1WDU3IIM+Ws8iLfYyWDzGaWks/2C5RVVYooAmFw7i
kXhJOGIeI5O7KB8vp//PndciBdymztME+E2K9rYGXRZrWOcU8wHCK432IU2C9kxk
Zt8k1KbhuSbjr0LACUdvo7ow64JjDtyBwoM9BRo9eTHFPqVkpGYvU+guqzM3uMzT
sXAiyCAIJeRVWSfqXG//M2G0D9dwTTtEhLq2PfBn5Tt2JGpAVOVLHY1wrWhoDmQq
sCU0kAWdjPXEJJB1UMK39uKIoXvVLPTCMom5U/dgEt4wkLO3hR9VtOv/3oW02wYw
lKrp9e2GsA0OOX2S0k2IAP0bYy9lR6rFX3TZPXPm/f+IMDxy8/J+CzUVRsHJvEcw
3dE7HQ8c3OQACyzG9wK6F7PYibfiA4qR3+u1BJWHmb9uXcmXL3jhxePWfidO3yMS
2AXduEe5gC6hYN+JQKyWDHgQ9oD3mCNbCZlJjQdIF/wFuBZ9zO02fmdBcGpCnacu
6moDLdtwHeIGlsLvopOyVbM8vFZHbMyrrb9Zz9uUzKCg/ftkT1fADTHJss+P4bmL
KwJvz2NcakOtUW8PvR73I8a1OmRpo8ewL32pUeNqBW06ctPg08gbBjWufCc0WlGw
bMAxcxx0AT0YT/mXunACYb5jdmYi0snCDD7GlAAHpFO5OqWTA3AJ7ip5Is7yvhtK
BkqewTh8F71g1B+WMcDfxQeLqgXyEtmNJr+fISBvwub5iFsDjYmd/hC++3R2MNLq
CZjGXx/amQyDrZeVgFvDK0PyvWALkENI6WkPn+11XiV7V7poz5ExjuEYGlVLGKlS
VrxxHobqOSbB/HLtTXsNexb4kYfQD14IO7zTAu5HrFzbl/rwiaWp2okjQwqhb/Gs
NLX2eSJZYIT2nmLH0o/mKEAz1IAx6tRJ+Gh/3X4LAoxIIzXcc03qe5+nzXij8J8Q
QVT5HtxWlulQpI75BOTRYloNCfstV6BZqL//s8b6EEebR2XuB7sKmoIWLl2M9UTg
fYTXSesh8bwee5Zzzc/6GdCS3VFOViJcGnaqdWGrDqp/b4jjmeIFwIAsRigBh8fC
rHO16js1DbTAAU0+fp+SS3SgKf3uEIMQ3dHVWFZPenI8zqTMoigQCJri3ydK1+Dt
rhaQJlRSscRQN95oEZr9/odk1xayWEJUP/2sxv3cKGWh9EIP8maAwhHgdcG4AnKO
+PUejOrEfLTMIDDCP4G4SqqS6CX7p9FrIvEy6FSk3TIShU7bs3MRW5rraR99iLwg
gvqSBKGgrqtZMxjRMKLOe5O65QpiqJmd9KQBUh6dVB2CTSpfhMDwB5wiCODtfqRx
zeuKx2MmcP8D0KGjIICX1ZIi46hrINXK96WfO1EO3O8CrNxEGNXdHJV9DT6mXRDk
Lw7sk909P7BMtZXyyOvq4hlZ2GaVmg1sACx4bLonEOMiS4d8EKFUVkpHDQXw0t1k
4rKPUu4EW77X/mCbqtcIqkKwfYZwSSlF8EnOJUTtr60v8jAuXnhMNSwiP/6hGxyB
/4N3QyMzAsPCBSoJ1srVK/kdY0PCioHn7PDcpIFo0MWegrXcWzX/fyTe1Q3D8Gkr
u2j4sCFaBxDRHttumd4VT0DNWUTZ1r871N6yN85W8kIj0HeRhj7PsYJAEfG6Jsdm
XrReUCch2HX11fB+RT6QgJiaPm/yoM9eI4gFlJb3iNJJPVzUGAgMOCVCRM4wAahV
zfCcIqvDjxWdYkAoJGRi+9UODl6BnOX32Db+hxNCIrS3kxZRf4MXG8dVRRlBIkPb
m6nKyY27bGazhttEmuKG06zl0dGUJkEnOdOxpy77yN1ys6+LY7w1zK1OvYB4G0ss
I6++ZTSeihMORcfKx0jyT4PjxYeXLpe9yrCaxhgylAgq2M8gO69uiAV/GrdBldkD
JgTXDsJCIyyideOAC5W1SX3OvEPUd76VcvLWCmU6+u/IVRXAQMc1f8+LKqetK+5T
b6hKpnPwRgJtftQbWwVlbMWL8p2FM36eJkH5uXfgCamssAE4AAp7O9ebxuZoSiLm
AaWpfpIKRbKWyYyufZWtvTnyVjDfApubcpiUTxl0qdeF8LmybBoGLe5xgDrOdBHM
CxWoR5105z1OX75kW8vmLQpgNrv+LTWJvgan/l8a6777jHVGbcskOaCRHw4NFKZg
zhDmFFFg1fORKGHpBWsGh0nERty/ehGASZwgY2lO+NM/p4OoGTp9RNoGQBict4/g
+CLxU0zXMuxjMxB50qsZXG7UY0UZ84tDUmCcEBAccAtB+L536pamY99ZYOB8Qi3+
bC1rJqo38JSyp+Qpv9OkDFgrSlMtgkFXiRMAEYB7J5xiGfZs4qebNoWVeIm68Ydt
s2dH8TRpM13AYwML2yWCv+XqXYOrjSfH/MF+zOiefslC/fMmZIseYJ98Z1NNa9pM
SBHwqwwJZe2p7tWJsImzBSWUMYljip/uYFY2aooeYV0OzdODiNEs3zED2tgvJUJ6
bgWR6pYQQo8BASYV6JNG1DhCqIP6TRV0Wg6vd6cKL/i7sozGo+Y5Ir8+G1Ynl1FV
WooucGkO5UyOx14oYsFWziSXCCVeBJZ8P7hysab0f0cw0kK9qXoJCCMha37T4YS6
TXr5vl/K845WNJn2FPmi0kF29vQ7yAHVWBux+hQ65EwdUR4eEsreuSkdA0yWScpi
TcsPuKBz3y2TzZbdcqeeCPG5KqThO60Y6CIrSg6o0ZN7kFQ32IaCogxLncapjKHh
p4NkvEuI7ZObQHz0XGVeEWxkFMangc0ud4iiBLQi1S35TZbVMZKuSOZ8wFQG+aZA
uWkQ1eX7ELyfGrVRB0cMP5OuK/2s5KfIC/+yS6/66OgsihIegncA0fn+veHexNId
3D0Kwcn8XPhWCuj3yD+YJg0ZsC8yJXSWIFOQWw8r9i5YBLd5Gr5p4/v2sSxgFzrg
JOMglL1RSredH/aUSc0T6vRhy83zcRwE5eXsYLXdFymxAGO5QhYcARtC+kIPHU94
Ze3npwHvELAg8e3s+JpM4DK+4BVkmQZXsKHULVXATnEMA69bVIvp6znLa9exFLbv
01wgai/Yz63B3BNWXt+/4n9LbpUHddvKAS00V42xee5/SJ2KoKH4RCzcSA3R1V/e
ql0iNoXOxmLCtNLtx/zxfwLM1ll6w1w7PgYqx0O6YctIK/iwx0GzLEEfMQmEB6E/
5pbrkVyW4G/KqU19HuifDnK+/pn7AvxOL0GQK5fy0UjrwHngssyCGHGnk9xVN8h3
+mSJfoaEsKa/Vps0xTTxqp+tKXGPV8In91mli5mEHNuXv8jn7mEmrGN0ATuiz2vU
BlXaON+bW55LciXTNtveknmiuK9NqKO7+xh2YLkjPOx1J3fag5a7kqtx22yyAC5h
6FIvfYU4oI2jOXJmzlLahvG7IpgfbfSpQOgU0SjgW3jJwMD2MNMirLkaBX4rrSq8
wukl1D2hYqhF+bPTEd1kLNbQYuYERx6runTT5C5eTzezTeFv/bMZwaC158oY7uLb
5oElKQaOjrwJsVunGEQnjAOggF9Lula5133BdPLaYwoTN6v9pZ2Kbx+nspBmJ4Vm
RJWVqVgljml1/b2xL1EGK9PxkNgvb91qefO0GPn6Nkr1A3TjsDwClz3ora3xcgOd
brvszTPMhT2Ay6gyVgOiZMzaxxX7jc96l5fBkJu6mONhDGppuorTGWQzLaxfDtT1
EWcRicSQWZb+/NLQqlOhqHQzD1zDqXqTGGhH7UrhKqGugd//+fIf3DYl9cX2b1BT
eYAR4i4pGI9xprottRwH2/6blH6aa6vR9xzyRp2aBLfjI01wEJ4oMdw3EHO43v5V
XAL0P+tS/ZJPOXxLMysrX+pg0mRG8fZxvtjaX82hKsbW0GSSX4YEnZ3QJzaC4Pdp
0Bx3HiiFWdE2dStrpbcoLiDnG8ONOeM660Oy/6feWmM49INbmK50L5y/G1tBQpV8
PpZPmgLZCgOwWVrBP+DhITAy7LzRsonty7NcROpbnALYj5Eyl8TV8+wXznW5tRHG
5KRavc3PtMDTsm7X7gouauH2SoJIz0G379cH9nagXeyuMlEFEeVqlt2AS2cvkp68
4H2xVwSrFAj+sTHbC07MT8ZnMo1rQ1oeq9IRB2aFGVxeJbfWab/sdgbM2Ou9y7b+
W6llTaW8p5FIJKa+EODpM9hREHtOzliWz3yyOsHsWxDk4QBkSiPn+swviKltaV//
BtbyBrcC3d4U5trCG1rgut3OpRUIyUosdZsIYFHlkLWZCQYmLApqjJgHusLuOjs8
IBubgSLJx+fJCWSW9VZ4aURc87aS8dLZwFoeXMaBv4ZiMoR+S9YzYw4EBju08MfE
v5lc5WF7vX3TQYeeiiMHO/ndu06q6mwAlOPxFe23uvaU8x7A4jJkirJQDaxc5FmL
hVWN7T6ERCZHUTstY8uQ1K18A0BpXqXPhhzZ484ImAQUhlHLrYKQ9Y8knU8fYxW8
EvRGHXUeKU1SRMXGkH2j2Bgz7XsEsYbMS6ucQVaycNNpg3Ebo5M/8+f3NB6DoDUV
S8RmbL4ggkK8RFfULtAGuIQJ/2wziKPIsEx8lgWAXsQQTlJrXyN/uPSuAVJHHD1+
wA3CP57S71b2xGpTImGLJ6dzjOEijD0+Ade0GYk5JaU/xZV+hgJidDENO5d+EZsY
VjM+iDiczUmz14yX+351EAjKkH/Zjn+dFziBNORwmP11+V6OYoDpgA3LKpEWvdIp
z3+FPhK0N108Oq5utFtMx1kggL6uu2vZms38JbSkIuWHiIsbkt7yQ1niHuBwROLp
57uINx6+D9dBVnVC5cw9LPeHVl7Z0WOaPnds13SJmlfllN473AKidQB1eJ/0fS/z
I1cZkd43brr8kvujFdTD3I57E/Zq+sMslqEclL5cxThhDdFzA+Qv7prZ/xBFPRu3
tygTHU7wC61RpV9EuToL8sKQwyL1eGjp0C4xCsNaSFkZ6vZpCVdADKgZCvWP1A5k
C65fJT1vNOQFlL66ycLcyoTJ9D+62fgjoivpQPGtwkSz/8svxSo3jcDWtSFKhm+m
9hSo7pQXoQwnX63UvcCg59RIPRNq/TLmCeVZdbbfUiEKvvsOTyiStEvoEkW5CG+P
+SwGDxmAlk/1nDXDWha6bG9WGSbw2BJ0Bz1bQ4o8eVkauRzUP/mBtrTy3QON/HVl
KsAxzMo89I2TCe7iIBsI4n+WaK3L1IhAAFStc+Fn0gvWb2QJ27dT2VH+5ilpVJkb
80rzicdTwGXHt6nNAxo7Z9da6vXWMYGo6GIolSKo0KZ+ReB1vOn8ryi/fiZAICPz
HmjcUYKr18QyRI0B6V2w93dBcbR9kXJdq/WoTgh4NseRYSF3b8cczyQfmn3lEAty
mNl4F/RrHXIIrWT7nQ1LBwZukYcGrjRog8C+dOjVJNN+APE2NsZo1QfycOioe8au
iHp7IL197Y2ePvj0rOJ8JjjetJCrKnTFzNnAlnfzqLhjKdzWjYXcGFUT/groFn4L
naP08q9ZlV6ZxTUWv5odJqv3g77id44MoR56qujf42Vlyh7U/5RZN57Ht89NJMjD
IHs+u2DsRcs6KxOdhtVvGmEGRWUYGUpQajb7rpbEMfvQhhrkqQFz0Uq9pUI2LmtD
o+E6QP+4kMSU8apuY4+BHr5ScsZA/MhvnWcR7QmQobsrr+1ojKTN0mCy+vLZhlEJ
f1nWrtdc+S3qDTeCBHGWoVeh0qKStDLHxikOORhjp8CzPR8KkQYdfPiuECrkCP//
LagOxfDhY2b1YWyPDsdjamCDgVYuP4T/kzt3gttZ7k6Dx8UbqVa4W6E+/hutKyZb
0MQWqxXG8BWavOAAtXK6eI+y0wyrO+uaNWufvguLjmm9/dXAwTWkJJzVaH2HVWVX
vmY4yu/QO/FXWZTsIiF/qazi9WD3jG4F5TZiGyiwemIB9fAHWMKcz8N37kifB8Bp
7QSinDWYBwV4LFirpd9KPX2JcHyeGzIPyEY9/k8Hynga+2XGet5+T1t3ugpfq9J+
zG6PE+xX+BRX5sfXJj5y/LEt3pGNr7ebnVfV2aWvA2aj5NNK8U3UfFomsv8pwdgM
y2E2vOagBs4hhR9lN7ylofzf0egjr/Hxqvvyr+s8i76xnvOzBkehs+qJFAd9gPAY
+DIH14qM6hBHubdfRaU/zfeBftQZDxt2pKYemu9/I/N3EV7BHfiqmVZt06NccKmV
Lplhs7SsfyD0hhJuNpDPGzamsbNtQ2aLk9sTbP9smVSWdhVDO0+S+B7dPD8pDp1v
/QPb5cyy8W+eI3/4Xpt1xPhFG5SgF+r4WwdsZUWYsfIzZBfb3HJRM8PAgHHakE1/
0+BVwo1Jo8WSw6MpP+7pjGCbGy9ajBThvOmNJR1iRlu/fSvD9w4sZ2COKHLI7gNn
+Gebju8P0QT+JNZfna7ZDHFgvSUDo8NnYOll3Fd4HHYt7gYd8IJ3U+ehcoww2HWk
jDppgTtFlNmb/NB3/f71q9GDX9vZ8mKiRXJYSYIhFTxGhBQMmtEPw5EUzr+7eolf
uf/D+VCpi0UWbiY0A7hKlM7Uq+pNQpYmtAU9rzfVCrOBV3x51JQqlcetFi8kmD1t
/rE4SW11cNWDwK13SMpAmibnpXGP20Tzg/6QQJOkZMyeqYd4MxfYl2EifxVwXHG6
aeW19rAwLqhJpIAU8GFp83d+9+dYJ3QLBAQhPgF+VE5KhhVkmESRw3oVtI5P1ckh
v8xr/2JCznTH0tG2/XwyzyK6IdVfBmMIvniPNg2RtKTG6VzMFJ3xWN+LUKvOAMw0
4CtzA2lXaoU0Fz+GLotOWh+WqAbJsdhDHJGS3v+YiWihiP8MlZ6z1JVwxlPs1yug
`pragma protect end_protected
